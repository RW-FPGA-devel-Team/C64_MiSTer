-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c5",
     9 => x"d4080b0b",
    10 => x"80c5d808",
    11 => x"0b0b80c5",
    12 => x"dc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c5dc0c0b",
    16 => x"0b80c5d8",
    17 => x"0c0b0b80",
    18 => x"c5d40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb498",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c5d470",
    57 => x"80d08427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5189dd",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c5",
    65 => x"e40c9f0b",
    66 => x"80c5e80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c5e808ff",
    70 => x"0580c5e8",
    71 => x"0c80c5e8",
    72 => x"088025e8",
    73 => x"3880c5e4",
    74 => x"08ff0580",
    75 => x"c5e40c80",
    76 => x"c5e40880",
    77 => x"25d03880",
    78 => x"0b80c5e8",
    79 => x"0c800b80",
    80 => x"c5e40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c5e408",
   100 => x"25913882",
   101 => x"c82d80c5",
   102 => x"e408ff05",
   103 => x"80c5e40c",
   104 => x"838a0480",
   105 => x"c5e40880",
   106 => x"c5e80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c5e408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c5e80881",
   116 => x"0580c5e8",
   117 => x"0c80c5e8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c5e8",
   121 => x"0c80c5e4",
   122 => x"08810580",
   123 => x"c5e40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c5",
   128 => x"e8088105",
   129 => x"80c5e80c",
   130 => x"80c5e808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c5e8",
   134 => x"0c80c5e4",
   135 => x"08810580",
   136 => x"c5e40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"c5ec0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"c5ec0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280c5",
   177 => x"ec088407",
   178 => x"80c5ec0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b0bbe",
   183 => x"9c0c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80c5ec",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80c5",
   208 => x"d40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050d84bf",
   216 => x"5186c72d",
   217 => x"ff115170",
   218 => x"8025f638",
   219 => x"0284050d",
   220 => x"0402fc05",
   221 => x"0dec5183",
   222 => x"710c86c7",
   223 => x"2d82710c",
   224 => x"909c2d02",
   225 => x"84050d04",
   226 => x"02fc050d",
   227 => x"ec518182",
   228 => x"710c86c7",
   229 => x"2d82710c",
   230 => x"909c2d02",
   231 => x"84050d04",
   232 => x"02fc050d",
   233 => x"ec5180c2",
   234 => x"710c86c7",
   235 => x"2d82710c",
   236 => x"909c2d02",
   237 => x"84050d04",
   238 => x"02fc050d",
   239 => x"ec518282",
   240 => x"710c86c7",
   241 => x"2d82710c",
   242 => x"909c2d02",
   243 => x"84050d04",
   244 => x"02fc050d",
   245 => x"ec519271",
   246 => x"0c86c72d",
   247 => x"82710c02",
   248 => x"84050d04",
   249 => x"02d0050d",
   250 => x"7d548074",
   251 => x"5380c5f0",
   252 => x"525bab82",
   253 => x"2d80c5d4",
   254 => x"087b2e81",
   255 => x"b63880c5",
   256 => x"f40870f8",
   257 => x"0c891580",
   258 => x"f52d8a16",
   259 => x"80f52d71",
   260 => x"82802905",
   261 => x"881780f5",
   262 => x"2d708480",
   263 => x"802912f4",
   264 => x"0c575556",
   265 => x"58a40bec",
   266 => x"0c7aff19",
   267 => x"585a767b",
   268 => x"2e8b3881",
   269 => x"1a77812a",
   270 => x"585a76f7",
   271 => x"38f71a5a",
   272 => x"815b8078",
   273 => x"2580ec38",
   274 => x"79527651",
   275 => x"84a82d80",
   276 => x"c6bc5280",
   277 => x"c5f051ad",
   278 => x"cf2d80c5",
   279 => x"d408802e",
   280 => x"b93880c6",
   281 => x"bc5c83fc",
   282 => x"597b7084",
   283 => x"055d0870",
   284 => x"81ff0671",
   285 => x"882a7081",
   286 => x"ff067390",
   287 => x"2a7081ff",
   288 => x"0675982a",
   289 => x"e80ce80c",
   290 => x"58e80c57",
   291 => x"e80cfc1a",
   292 => x"5a537880",
   293 => x"25d33889",
   294 => x"a20480c5",
   295 => x"d4085b84",
   296 => x"805880c5",
   297 => x"f051ad9f",
   298 => x"2dfc8018",
   299 => x"81185858",
   300 => x"88c20486",
   301 => x"da2d840b",
   302 => x"ec0c7a80",
   303 => x"2e8e3880",
   304 => x"c1c45192",
   305 => x"a62d909c",
   306 => x"2d89d304",
   307 => x"80c3a451",
   308 => x"92a62d7a",
   309 => x"80c5d40c",
   310 => x"02b0050d",
   311 => x"0402ec05",
   312 => x"0d840bec",
   313 => x"0c8ffa2d",
   314 => x"8ccc2d81",
   315 => x"f92da1c2",
   316 => x"2d80c5d4",
   317 => x"08802e82",
   318 => x"bc3887e4",
   319 => x"51b48f2d",
   320 => x"80c1c451",
   321 => x"92a62d90",
   322 => x"9c2d8cd8",
   323 => x"2d92b92d",
   324 => x"80c0b80b",
   325 => x"80f52d70",
   326 => x"822b8406",
   327 => x"80c0c40b",
   328 => x"80f52d70",
   329 => x"982b8180",
   330 => x"0a0680c0",
   331 => x"d00b80f5",
   332 => x"2d70842b",
   333 => x"b0067473",
   334 => x"070780c0",
   335 => x"dc0b80f5",
   336 => x"2d70882b",
   337 => x"86800680",
   338 => x"c0e80b80",
   339 => x"f52d7372",
   340 => x"07719e2b",
   341 => x"07bf980b",
   342 => x"80f52d70",
   343 => x"8d2b80c0",
   344 => x"8006bfa4",
   345 => x"0b80f52d",
   346 => x"70902b84",
   347 => x"80800674",
   348 => x"730707bf",
   349 => x"b00b80f5",
   350 => x"2d70942b",
   351 => x"98800a06",
   352 => x"bfbc0b80",
   353 => x"f52d708c",
   354 => x"2ba08006",
   355 => x"74730707",
   356 => x"bfc80b80",
   357 => x"f52d7092",
   358 => x"2bb08080",
   359 => x"06bfd40b",
   360 => x"80f52d70",
   361 => x"962b8680",
   362 => x"0a067473",
   363 => x"0707bea8",
   364 => x"0b80f52d",
   365 => x"70832b88",
   366 => x"06beb40b",
   367 => x"80f52d70",
   368 => x"10820674",
   369 => x"730707be",
   370 => x"c00b80f5",
   371 => x"2d709a2b",
   372 => x"b00a06be",
   373 => x"cc0b80f5",
   374 => x"2d709c2b",
   375 => x"8c0a0674",
   376 => x"73070780",
   377 => x"c2ac0b80",
   378 => x"f52d708e",
   379 => x"2b838080",
   380 => x"0680c2b8",
   381 => x"0b80f52d",
   382 => x"708b2b90",
   383 => x"80067473",
   384 => x"0707fc0c",
   385 => x"54545454",
   386 => x"54545454",
   387 => x"54545454",
   388 => x"54545454",
   389 => x"54545454",
   390 => x"54555354",
   391 => x"54575354",
   392 => x"52575753",
   393 => x"53865280",
   394 => x"c5d40883",
   395 => x"38845271",
   396 => x"ec0c8a8a",
   397 => x"04800b80",
   398 => x"c5d40c02",
   399 => x"94050d04",
   400 => x"71980c04",
   401 => x"ffb00880",
   402 => x"c5d40c04",
   403 => x"810bffb0",
   404 => x"0c04800b",
   405 => x"ffb00c04",
   406 => x"02f4050d",
   407 => x"8de60480",
   408 => x"c5d40881",
   409 => x"f02e0981",
   410 => x"068a3881",
   411 => x"0b80c488",
   412 => x"0c8de604",
   413 => x"80c5d408",
   414 => x"81e02e09",
   415 => x"81068a38",
   416 => x"810b80c4",
   417 => x"8c0c8de6",
   418 => x"0480c5d4",
   419 => x"085280c4",
   420 => x"8c08802e",
   421 => x"893880c5",
   422 => x"d4088180",
   423 => x"05527184",
   424 => x"2c728f06",
   425 => x"535380c4",
   426 => x"8808802e",
   427 => x"9a387284",
   428 => x"2980c3c8",
   429 => x"05721381",
   430 => x"712b7009",
   431 => x"73080673",
   432 => x"0c515353",
   433 => x"8dda0472",
   434 => x"842980c3",
   435 => x"c8057213",
   436 => x"83712b72",
   437 => x"0807720c",
   438 => x"5353800b",
   439 => x"80c48c0c",
   440 => x"800b80c4",
   441 => x"880c80c5",
   442 => x"fc518eed",
   443 => x"2d80c5d4",
   444 => x"08ff24fe",
   445 => x"ea38800b",
   446 => x"80c5d40c",
   447 => x"028c050d",
   448 => x"0402f805",
   449 => x"0d80c3c8",
   450 => x"528f5180",
   451 => x"72708405",
   452 => x"540cff11",
   453 => x"51708025",
   454 => x"f2380288",
   455 => x"050d0402",
   456 => x"f0050d75",
   457 => x"518cd22d",
   458 => x"70822cfc",
   459 => x"0680c3c8",
   460 => x"1172109e",
   461 => x"06710870",
   462 => x"722a7083",
   463 => x"0682742b",
   464 => x"70097406",
   465 => x"760c5451",
   466 => x"56575351",
   467 => x"538ccc2d",
   468 => x"7180c5d4",
   469 => x"0c029005",
   470 => x"0d0402fc",
   471 => x"050d7251",
   472 => x"80710c80",
   473 => x"0b84120c",
   474 => x"0284050d",
   475 => x"0402f005",
   476 => x"0d757008",
   477 => x"84120853",
   478 => x"5353ff54",
   479 => x"71712ea8",
   480 => x"388cd22d",
   481 => x"84130870",
   482 => x"84291488",
   483 => x"11700870",
   484 => x"81ff0684",
   485 => x"18088111",
   486 => x"8706841a",
   487 => x"0c535155",
   488 => x"5151518c",
   489 => x"cc2d7154",
   490 => x"7380c5d4",
   491 => x"0c029005",
   492 => x"0d0402f8",
   493 => x"050d8cd2",
   494 => x"2de00870",
   495 => x"8b2a7081",
   496 => x"06515252",
   497 => x"70802ea1",
   498 => x"3880c5fc",
   499 => x"08708429",
   500 => x"80c68405",
   501 => x"7381ff06",
   502 => x"710c5151",
   503 => x"80c5fc08",
   504 => x"81118706",
   505 => x"80c5fc0c",
   506 => x"51800b80",
   507 => x"c6a40c8c",
   508 => x"c42d8ccc",
   509 => x"2d028805",
   510 => x"0d0402fc",
   511 => x"050d80c5",
   512 => x"fc518eda",
   513 => x"2d8e812d",
   514 => x"8fb2518c",
   515 => x"c02d0284",
   516 => x"050d0480",
   517 => x"c6a80880",
   518 => x"c5d40c04",
   519 => x"02fc050d",
   520 => x"90a6048c",
   521 => x"d82d80f6",
   522 => x"518e9f2d",
   523 => x"80c5d408",
   524 => x"f23880da",
   525 => x"518e9f2d",
   526 => x"80c5d408",
   527 => x"e63880c5",
   528 => x"d40880c4",
   529 => x"940c80c5",
   530 => x"d4085185",
   531 => x"8d2d0284",
   532 => x"050d0402",
   533 => x"ec050d76",
   534 => x"54805287",
   535 => x"0b881580",
   536 => x"f52d5653",
   537 => x"74722483",
   538 => x"38a05372",
   539 => x"5183842d",
   540 => x"81128b15",
   541 => x"80f52d54",
   542 => x"52727225",
   543 => x"de380294",
   544 => x"050d0402",
   545 => x"f0050d80",
   546 => x"c6a80854",
   547 => x"81f92d80",
   548 => x"0b80c6ac",
   549 => x"0c730880",
   550 => x"2e818638",
   551 => x"820b80c5",
   552 => x"e80c80c6",
   553 => x"ac088f06",
   554 => x"80c5e40c",
   555 => x"73085271",
   556 => x"832e9638",
   557 => x"71832689",
   558 => x"3871812e",
   559 => x"af38928a",
   560 => x"0471852e",
   561 => x"9f38928a",
   562 => x"04881480",
   563 => x"f52d8415",
   564 => x"08bce853",
   565 => x"545286a0",
   566 => x"2d718429",
   567 => x"13700852",
   568 => x"52928e04",
   569 => x"735190d3",
   570 => x"2d928a04",
   571 => x"80c49008",
   572 => x"8815082c",
   573 => x"70810651",
   574 => x"5271802e",
   575 => x"8738bcec",
   576 => x"51928704",
   577 => x"bcf05186",
   578 => x"a02d8414",
   579 => x"085186a0",
   580 => x"2d80c6ac",
   581 => x"08810580",
   582 => x"c6ac0c8c",
   583 => x"14549195",
   584 => x"04029005",
   585 => x"0d047180",
   586 => x"c6a80c91",
   587 => x"832d80c6",
   588 => x"ac08ff05",
   589 => x"80c6b00c",
   590 => x"0402e805",
   591 => x"0d80c6a8",
   592 => x"0880c6b4",
   593 => x"08575587",
   594 => x"518e9f2d",
   595 => x"80c5d408",
   596 => x"812a7081",
   597 => x"06515271",
   598 => x"802ea338",
   599 => x"92e2048c",
   600 => x"d82d8751",
   601 => x"8e9f2d80",
   602 => x"c5d408f3",
   603 => x"3880c494",
   604 => x"08813270",
   605 => x"80c4940c",
   606 => x"70525285",
   607 => x"8d2d80fe",
   608 => x"518e9f2d",
   609 => x"80c5d408",
   610 => x"802ea938",
   611 => x"80c49408",
   612 => x"802e9238",
   613 => x"800b80c4",
   614 => x"940c8051",
   615 => x"858d2d93",
   616 => x"a5048cd8",
   617 => x"2d80fe51",
   618 => x"8e9f2d80",
   619 => x"c5d408f2",
   620 => x"3887d02d",
   621 => x"80c49408",
   622 => x"903881fd",
   623 => x"518e9f2d",
   624 => x"81fa518e",
   625 => x"9f2d999e",
   626 => x"0481f551",
   627 => x"8e9f2d80",
   628 => x"c5d40881",
   629 => x"2a708106",
   630 => x"51527180",
   631 => x"2eb33880",
   632 => x"c6b00852",
   633 => x"71802e8a",
   634 => x"38ff1280",
   635 => x"c6b00c94",
   636 => x"910480c6",
   637 => x"ac081080",
   638 => x"c6ac0805",
   639 => x"70842916",
   640 => x"51528812",
   641 => x"08802e89",
   642 => x"38ff5188",
   643 => x"12085271",
   644 => x"2d81f251",
   645 => x"8e9f2d80",
   646 => x"c5d40881",
   647 => x"2a708106",
   648 => x"51527180",
   649 => x"2eb43880",
   650 => x"c6ac08ff",
   651 => x"1180c6b0",
   652 => x"08565353",
   653 => x"7372258a",
   654 => x"38811480",
   655 => x"c6b00c94",
   656 => x"da047210",
   657 => x"13708429",
   658 => x"16515288",
   659 => x"1208802e",
   660 => x"8938fe51",
   661 => x"88120852",
   662 => x"712d81fd",
   663 => x"518e9f2d",
   664 => x"80c5d408",
   665 => x"812a7081",
   666 => x"06515271",
   667 => x"802eb138",
   668 => x"80c6b008",
   669 => x"802e8a38",
   670 => x"800b80c6",
   671 => x"b00c95a0",
   672 => x"0480c6ac",
   673 => x"081080c6",
   674 => x"ac080570",
   675 => x"84291651",
   676 => x"52881208",
   677 => x"802e8938",
   678 => x"fd518812",
   679 => x"0852712d",
   680 => x"81fa518e",
   681 => x"9f2d80c5",
   682 => x"d408812a",
   683 => x"70810651",
   684 => x"5271802e",
   685 => x"b13880c6",
   686 => x"ac08ff11",
   687 => x"545280c6",
   688 => x"b0087325",
   689 => x"89387280",
   690 => x"c6b00c95",
   691 => x"e6047110",
   692 => x"12708429",
   693 => x"16515288",
   694 => x"1208802e",
   695 => x"8938fc51",
   696 => x"88120852",
   697 => x"712d80c6",
   698 => x"b0087053",
   699 => x"5473802e",
   700 => x"8a388c15",
   701 => x"ff155555",
   702 => x"95ed0482",
   703 => x"0b80c5e8",
   704 => x"0c718f06",
   705 => x"80c5e40c",
   706 => x"81eb518e",
   707 => x"9f2d80c5",
   708 => x"d408812a",
   709 => x"70810651",
   710 => x"5271802e",
   711 => x"ad387408",
   712 => x"852e0981",
   713 => x"06a43888",
   714 => x"1580f52d",
   715 => x"ff055271",
   716 => x"881681b7",
   717 => x"2d71982b",
   718 => x"52718025",
   719 => x"8838800b",
   720 => x"881681b7",
   721 => x"2d745190",
   722 => x"d32d81f4",
   723 => x"518e9f2d",
   724 => x"80c5d408",
   725 => x"812a7081",
   726 => x"06515271",
   727 => x"802eb338",
   728 => x"7408852e",
   729 => x"098106aa",
   730 => x"38881580",
   731 => x"f52d8105",
   732 => x"52718816",
   733 => x"81b72d71",
   734 => x"81ff068b",
   735 => x"1680f52d",
   736 => x"54527272",
   737 => x"27873872",
   738 => x"881681b7",
   739 => x"2d745190",
   740 => x"d32d80da",
   741 => x"518e9f2d",
   742 => x"80c5d408",
   743 => x"812a7081",
   744 => x"06515271",
   745 => x"802e81ad",
   746 => x"3880c6a8",
   747 => x"0880c6b0",
   748 => x"08555373",
   749 => x"802e8a38",
   750 => x"8c13ff15",
   751 => x"555397b3",
   752 => x"04720852",
   753 => x"71822ea6",
   754 => x"38718226",
   755 => x"89387181",
   756 => x"2eaa3898",
   757 => x"d5047183",
   758 => x"2eb43871",
   759 => x"842e0981",
   760 => x"0680f238",
   761 => x"88130851",
   762 => x"92a62d98",
   763 => x"d50480c6",
   764 => x"b0085188",
   765 => x"13085271",
   766 => x"2d98d504",
   767 => x"810b8814",
   768 => x"082b80c4",
   769 => x"90083280",
   770 => x"c4900c98",
   771 => x"a9048813",
   772 => x"80f52d81",
   773 => x"058b1480",
   774 => x"f52d5354",
   775 => x"71742483",
   776 => x"38805473",
   777 => x"881481b7",
   778 => x"2d91832d",
   779 => x"98d50475",
   780 => x"08802ea4",
   781 => x"38750851",
   782 => x"8e9f2d80",
   783 => x"c5d40881",
   784 => x"06527180",
   785 => x"2e8c3880",
   786 => x"c6b00851",
   787 => x"84160852",
   788 => x"712d8816",
   789 => x"5675d838",
   790 => x"8054800b",
   791 => x"80c5e80c",
   792 => x"738f0680",
   793 => x"c5e40ca0",
   794 => x"527380c6",
   795 => x"b0082e09",
   796 => x"81069938",
   797 => x"80c6ac08",
   798 => x"ff057432",
   799 => x"70098105",
   800 => x"7072079f",
   801 => x"2a917131",
   802 => x"51515353",
   803 => x"71518384",
   804 => x"2d811454",
   805 => x"8e7425c2",
   806 => x"3880c494",
   807 => x"08527180",
   808 => x"c5d40c02",
   809 => x"98050d04",
   810 => x"02f4050d",
   811 => x"d45281ff",
   812 => x"720c7108",
   813 => x"5381ff72",
   814 => x"0c72882b",
   815 => x"83fe8006",
   816 => x"72087081",
   817 => x"ff065152",
   818 => x"5381ff72",
   819 => x"0c727107",
   820 => x"882b7208",
   821 => x"7081ff06",
   822 => x"51525381",
   823 => x"ff720c72",
   824 => x"7107882b",
   825 => x"72087081",
   826 => x"ff067207",
   827 => x"80c5d40c",
   828 => x"5253028c",
   829 => x"050d0402",
   830 => x"f4050d74",
   831 => x"767181ff",
   832 => x"06d40c53",
   833 => x"5380c6b8",
   834 => x"08853871",
   835 => x"892b5271",
   836 => x"982ad40c",
   837 => x"71902a70",
   838 => x"81ff06d4",
   839 => x"0c517188",
   840 => x"2a7081ff",
   841 => x"06d40c51",
   842 => x"7181ff06",
   843 => x"d40c7290",
   844 => x"2a7081ff",
   845 => x"06d40c51",
   846 => x"d4087081",
   847 => x"ff065151",
   848 => x"82b8bf52",
   849 => x"7081ff2e",
   850 => x"09810694",
   851 => x"3881ff0b",
   852 => x"d40cd408",
   853 => x"7081ff06",
   854 => x"ff145451",
   855 => x"5171e538",
   856 => x"7080c5d4",
   857 => x"0c028c05",
   858 => x"0d0402fc",
   859 => x"050d81c7",
   860 => x"5181ff0b",
   861 => x"d40cff11",
   862 => x"51708025",
   863 => x"f4380284",
   864 => x"050d0402",
   865 => x"f4050d81",
   866 => x"ff0bd40c",
   867 => x"93538052",
   868 => x"87fc80c1",
   869 => x"5199f72d",
   870 => x"80c5d408",
   871 => x"8b3881ff",
   872 => x"0bd40c81",
   873 => x"539bb104",
   874 => x"9aea2dff",
   875 => x"135372de",
   876 => x"387280c5",
   877 => x"d40c028c",
   878 => x"050d0402",
   879 => x"ec050d81",
   880 => x"0b80c6b8",
   881 => x"0c8454d0",
   882 => x"08708f2a",
   883 => x"70810651",
   884 => x"515372f3",
   885 => x"3872d00c",
   886 => x"9aea2dbc",
   887 => x"f45186a0",
   888 => x"2dd00870",
   889 => x"8f2a7081",
   890 => x"06515153",
   891 => x"72f33881",
   892 => x"0bd00cb1",
   893 => x"53805284",
   894 => x"d480c051",
   895 => x"99f72d80",
   896 => x"c5d40881",
   897 => x"2e933872",
   898 => x"822ebf38",
   899 => x"ff135372",
   900 => x"e438ff14",
   901 => x"5473ffaf",
   902 => x"389aea2d",
   903 => x"83aa5284",
   904 => x"9c80c851",
   905 => x"99f72d80",
   906 => x"c5d40881",
   907 => x"2e098106",
   908 => x"933899a8",
   909 => x"2d80c5d4",
   910 => x"0883ffff",
   911 => x"06537283",
   912 => x"aa2e9d38",
   913 => x"9b832d9c",
   914 => x"db04bd80",
   915 => x"5186a02d",
   916 => x"80539eb0",
   917 => x"04bd9851",
   918 => x"86a02d80",
   919 => x"549e8104",
   920 => x"81ff0bd4",
   921 => x"0cb1549a",
   922 => x"ea2d8fcf",
   923 => x"53805287",
   924 => x"fc80f751",
   925 => x"99f72d80",
   926 => x"c5d40855",
   927 => x"80c5d408",
   928 => x"812e0981",
   929 => x"069c3881",
   930 => x"ff0bd40c",
   931 => x"820a5284",
   932 => x"9c80e951",
   933 => x"99f72d80",
   934 => x"c5d40880",
   935 => x"2e8d389a",
   936 => x"ea2dff13",
   937 => x"5372c638",
   938 => x"9df40481",
   939 => x"ff0bd40c",
   940 => x"80c5d408",
   941 => x"5287fc80",
   942 => x"fa5199f7",
   943 => x"2d80c5d4",
   944 => x"08b23881",
   945 => x"ff0bd40c",
   946 => x"d4085381",
   947 => x"ff0bd40c",
   948 => x"81ff0bd4",
   949 => x"0c81ff0b",
   950 => x"d40c81ff",
   951 => x"0bd40c72",
   952 => x"862a7081",
   953 => x"06765651",
   954 => x"53729638",
   955 => x"80c5d408",
   956 => x"549e8104",
   957 => x"73822efe",
   958 => x"dc38ff14",
   959 => x"5473fee7",
   960 => x"387380c6",
   961 => x"b80c738b",
   962 => x"38815287",
   963 => x"fc80d051",
   964 => x"99f72d81",
   965 => x"ff0bd40c",
   966 => x"d008708f",
   967 => x"2a708106",
   968 => x"51515372",
   969 => x"f33872d0",
   970 => x"0c81ff0b",
   971 => x"d40c8153",
   972 => x"7280c5d4",
   973 => x"0c029405",
   974 => x"0d0402e8",
   975 => x"050d7855",
   976 => x"805681ff",
   977 => x"0bd40cd0",
   978 => x"08708f2a",
   979 => x"70810651",
   980 => x"515372f3",
   981 => x"3882810b",
   982 => x"d00c81ff",
   983 => x"0bd40c77",
   984 => x"5287fc80",
   985 => x"d15199f7",
   986 => x"2d80dbc6",
   987 => x"df5480c5",
   988 => x"d408802e",
   989 => x"8a38bdb8",
   990 => x"5186a02d",
   991 => x"9fd30481",
   992 => x"ff0bd40c",
   993 => x"d4087081",
   994 => x"ff065153",
   995 => x"7281fe2e",
   996 => x"0981069e",
   997 => x"3880ff53",
   998 => x"99a82d80",
   999 => x"c5d40875",
  1000 => x"70840557",
  1001 => x"0cff1353",
  1002 => x"728025ec",
  1003 => x"3881569f",
  1004 => x"b804ff14",
  1005 => x"5473c838",
  1006 => x"81ff0bd4",
  1007 => x"0c81ff0b",
  1008 => x"d40cd008",
  1009 => x"708f2a70",
  1010 => x"81065151",
  1011 => x"5372f338",
  1012 => x"72d00c75",
  1013 => x"80c5d40c",
  1014 => x"0298050d",
  1015 => x"0402e805",
  1016 => x"0d77797b",
  1017 => x"58555580",
  1018 => x"53727625",
  1019 => x"a3387470",
  1020 => x"81055680",
  1021 => x"f52d7470",
  1022 => x"81055680",
  1023 => x"f52d5252",
  1024 => x"71712e86",
  1025 => x"388151a0",
  1026 => x"92048113",
  1027 => x"539fe904",
  1028 => x"80517080",
  1029 => x"c5d40c02",
  1030 => x"98050d04",
  1031 => x"02ec050d",
  1032 => x"76557480",
  1033 => x"2e80c238",
  1034 => x"9a1580e0",
  1035 => x"2d51aea9",
  1036 => x"2d80c5d4",
  1037 => x"0880c5d4",
  1038 => x"0880ccec",
  1039 => x"0c80c5d4",
  1040 => x"08545480",
  1041 => x"ccc80880",
  1042 => x"2e9a3894",
  1043 => x"1580e02d",
  1044 => x"51aea92d",
  1045 => x"80c5d408",
  1046 => x"902b83ff",
  1047 => x"f00a0670",
  1048 => x"75075153",
  1049 => x"7280ccec",
  1050 => x"0c80ccec",
  1051 => x"08537280",
  1052 => x"2e9d3880",
  1053 => x"ccc008fe",
  1054 => x"14712980",
  1055 => x"ccd40805",
  1056 => x"80ccf00c",
  1057 => x"70842b80",
  1058 => x"cccc0c54",
  1059 => x"a1bd0480",
  1060 => x"ccd80880",
  1061 => x"ccec0c80",
  1062 => x"ccdc0880",
  1063 => x"ccf00c80",
  1064 => x"ccc80880",
  1065 => x"2e8b3880",
  1066 => x"ccc00884",
  1067 => x"2b53a1b8",
  1068 => x"0480cce0",
  1069 => x"08842b53",
  1070 => x"7280cccc",
  1071 => x"0c029405",
  1072 => x"0d0402d8",
  1073 => x"050d800b",
  1074 => x"80ccc80c",
  1075 => x"84549bbb",
  1076 => x"2d80c5d4",
  1077 => x"08802e97",
  1078 => x"3880c6bc",
  1079 => x"5280519e",
  1080 => x"ba2d80c5",
  1081 => x"d408802e",
  1082 => x"8638fe54",
  1083 => x"a1f704ff",
  1084 => x"14547380",
  1085 => x"24d83873",
  1086 => x"8c38bdc8",
  1087 => x"5186a02d",
  1088 => x"7355a7c4",
  1089 => x"04805681",
  1090 => x"0b80ccf4",
  1091 => x"0c8853bd",
  1092 => x"dc5280c6",
  1093 => x"f2519fdd",
  1094 => x"2d80c5d4",
  1095 => x"08762e09",
  1096 => x"81068938",
  1097 => x"80c5d408",
  1098 => x"80ccf40c",
  1099 => x"8853bde8",
  1100 => x"5280c78e",
  1101 => x"519fdd2d",
  1102 => x"80c5d408",
  1103 => x"893880c5",
  1104 => x"d40880cc",
  1105 => x"f40c80cc",
  1106 => x"f408802e",
  1107 => x"81803880",
  1108 => x"ca820b80",
  1109 => x"f52d80ca",
  1110 => x"830b80f5",
  1111 => x"2d71982b",
  1112 => x"71902b07",
  1113 => x"80ca840b",
  1114 => x"80f52d70",
  1115 => x"882b7207",
  1116 => x"80ca850b",
  1117 => x"80f52d71",
  1118 => x"0780caba",
  1119 => x"0b80f52d",
  1120 => x"80cabb0b",
  1121 => x"80f52d71",
  1122 => x"882b0753",
  1123 => x"5f54525a",
  1124 => x"56575573",
  1125 => x"81abaa2e",
  1126 => x"0981068e",
  1127 => x"387551ad",
  1128 => x"f82d80c5",
  1129 => x"d40856a3",
  1130 => x"b7047382",
  1131 => x"d4d52e87",
  1132 => x"38bdf451",
  1133 => x"a4800480",
  1134 => x"c6bc5275",
  1135 => x"519eba2d",
  1136 => x"80c5d408",
  1137 => x"5580c5d4",
  1138 => x"08802e83",
  1139 => x"f7388853",
  1140 => x"bde85280",
  1141 => x"c78e519f",
  1142 => x"dd2d80c5",
  1143 => x"d4088a38",
  1144 => x"810b80cc",
  1145 => x"c80ca486",
  1146 => x"048853bd",
  1147 => x"dc5280c6",
  1148 => x"f2519fdd",
  1149 => x"2d80c5d4",
  1150 => x"08802e8a",
  1151 => x"38be8851",
  1152 => x"86a02da4",
  1153 => x"e50480ca",
  1154 => x"ba0b80f5",
  1155 => x"2d547380",
  1156 => x"d52e0981",
  1157 => x"0680ce38",
  1158 => x"80cabb0b",
  1159 => x"80f52d54",
  1160 => x"7381aa2e",
  1161 => x"098106bd",
  1162 => x"38800b80",
  1163 => x"c6bc0b80",
  1164 => x"f52d5654",
  1165 => x"7481e92e",
  1166 => x"83388154",
  1167 => x"7481eb2e",
  1168 => x"8c388055",
  1169 => x"73752e09",
  1170 => x"810682f8",
  1171 => x"3880c6c7",
  1172 => x"0b80f52d",
  1173 => x"55748e38",
  1174 => x"80c6c80b",
  1175 => x"80f52d54",
  1176 => x"73822e86",
  1177 => x"388055a7",
  1178 => x"c40480c6",
  1179 => x"c90b80f5",
  1180 => x"2d7080cc",
  1181 => x"c00cff05",
  1182 => x"80ccc40c",
  1183 => x"80c6ca0b",
  1184 => x"80f52d80",
  1185 => x"c6cb0b80",
  1186 => x"f52d5876",
  1187 => x"05778280",
  1188 => x"29057080",
  1189 => x"ccd00c80",
  1190 => x"c6cc0b80",
  1191 => x"f52d7080",
  1192 => x"cce40c80",
  1193 => x"ccc80859",
  1194 => x"57587680",
  1195 => x"2e81b638",
  1196 => x"8853bde8",
  1197 => x"5280c78e",
  1198 => x"519fdd2d",
  1199 => x"80c5d408",
  1200 => x"82823880",
  1201 => x"ccc00870",
  1202 => x"842b80cc",
  1203 => x"cc0c7080",
  1204 => x"cce00c80",
  1205 => x"c6e10b80",
  1206 => x"f52d80c6",
  1207 => x"e00b80f5",
  1208 => x"2d718280",
  1209 => x"290580c6",
  1210 => x"e20b80f5",
  1211 => x"2d708480",
  1212 => x"80291280",
  1213 => x"c6e30b80",
  1214 => x"f52d7081",
  1215 => x"800a2912",
  1216 => x"7080cce8",
  1217 => x"0c80cce4",
  1218 => x"08712980",
  1219 => x"ccd00805",
  1220 => x"7080ccd4",
  1221 => x"0c80c6e9",
  1222 => x"0b80f52d",
  1223 => x"80c6e80b",
  1224 => x"80f52d71",
  1225 => x"82802905",
  1226 => x"80c6ea0b",
  1227 => x"80f52d70",
  1228 => x"84808029",
  1229 => x"1280c6eb",
  1230 => x"0b80f52d",
  1231 => x"70982b81",
  1232 => x"f00a0672",
  1233 => x"057080cc",
  1234 => x"d80cfe11",
  1235 => x"7e297705",
  1236 => x"80ccdc0c",
  1237 => x"52595243",
  1238 => x"545e5152",
  1239 => x"59525d57",
  1240 => x"5957a7bd",
  1241 => x"0480c6ce",
  1242 => x"0b80f52d",
  1243 => x"80c6cd0b",
  1244 => x"80f52d71",
  1245 => x"82802905",
  1246 => x"7080cccc",
  1247 => x"0c70a029",
  1248 => x"83ff0570",
  1249 => x"892a7080",
  1250 => x"cce00c80",
  1251 => x"c6d30b80",
  1252 => x"f52d80c6",
  1253 => x"d20b80f5",
  1254 => x"2d718280",
  1255 => x"29057080",
  1256 => x"cce80c7b",
  1257 => x"71291e70",
  1258 => x"80ccdc0c",
  1259 => x"7d80ccd8",
  1260 => x"0c730580",
  1261 => x"ccd40c55",
  1262 => x"5e515155",
  1263 => x"558051a0",
  1264 => x"9c2d8155",
  1265 => x"7480c5d4",
  1266 => x"0c02a805",
  1267 => x"0d0402ec",
  1268 => x"050d7670",
  1269 => x"872c7180",
  1270 => x"ff065556",
  1271 => x"5480ccc8",
  1272 => x"088a3873",
  1273 => x"882c7481",
  1274 => x"ff065455",
  1275 => x"80c6bc52",
  1276 => x"80ccd008",
  1277 => x"15519eba",
  1278 => x"2d80c5d4",
  1279 => x"085480c5",
  1280 => x"d408802e",
  1281 => x"b83880cc",
  1282 => x"c808802e",
  1283 => x"9a387284",
  1284 => x"2980c6bc",
  1285 => x"05700852",
  1286 => x"53adf82d",
  1287 => x"80c5d408",
  1288 => x"f00a0653",
  1289 => x"a8bb0472",
  1290 => x"1080c6bc",
  1291 => x"057080e0",
  1292 => x"2d5253ae",
  1293 => x"a92d80c5",
  1294 => x"d4085372",
  1295 => x"547380c5",
  1296 => x"d40c0294",
  1297 => x"050d0402",
  1298 => x"e0050d79",
  1299 => x"70842c80",
  1300 => x"ccf00805",
  1301 => x"718f0652",
  1302 => x"5553728a",
  1303 => x"3880c6bc",
  1304 => x"5273519e",
  1305 => x"ba2d72a0",
  1306 => x"2980c6bc",
  1307 => x"05548074",
  1308 => x"80f52d56",
  1309 => x"5374732e",
  1310 => x"83388153",
  1311 => x"7481e52e",
  1312 => x"81f43881",
  1313 => x"70740654",
  1314 => x"5872802e",
  1315 => x"81e8388b",
  1316 => x"1480f52d",
  1317 => x"70832a79",
  1318 => x"06585676",
  1319 => x"9b3880c4",
  1320 => x"98085372",
  1321 => x"89387280",
  1322 => x"cabc0b81",
  1323 => x"b72d7680",
  1324 => x"c4980c73",
  1325 => x"53aaf804",
  1326 => x"758f2e09",
  1327 => x"810681b6",
  1328 => x"38749f06",
  1329 => x"8d2980ca",
  1330 => x"af115153",
  1331 => x"811480f5",
  1332 => x"2d737081",
  1333 => x"055581b7",
  1334 => x"2d831480",
  1335 => x"f52d7370",
  1336 => x"81055581",
  1337 => x"b72d8514",
  1338 => x"80f52d73",
  1339 => x"70810555",
  1340 => x"81b72d87",
  1341 => x"1480f52d",
  1342 => x"73708105",
  1343 => x"5581b72d",
  1344 => x"891480f5",
  1345 => x"2d737081",
  1346 => x"055581b7",
  1347 => x"2d8e1480",
  1348 => x"f52d7370",
  1349 => x"81055581",
  1350 => x"b72d9014",
  1351 => x"80f52d73",
  1352 => x"70810555",
  1353 => x"81b72d92",
  1354 => x"1480f52d",
  1355 => x"73708105",
  1356 => x"5581b72d",
  1357 => x"941480f5",
  1358 => x"2d737081",
  1359 => x"055581b7",
  1360 => x"2d961480",
  1361 => x"f52d7370",
  1362 => x"81055581",
  1363 => x"b72d9814",
  1364 => x"80f52d73",
  1365 => x"70810555",
  1366 => x"81b72d9c",
  1367 => x"1480f52d",
  1368 => x"73708105",
  1369 => x"5581b72d",
  1370 => x"9e1480f5",
  1371 => x"2d7381b7",
  1372 => x"2d7780c4",
  1373 => x"980c8053",
  1374 => x"7280c5d4",
  1375 => x"0c02a005",
  1376 => x"0d0402cc",
  1377 => x"050d7e60",
  1378 => x"5e5a800b",
  1379 => x"80ccec08",
  1380 => x"80ccf008",
  1381 => x"595c5680",
  1382 => x"5880cccc",
  1383 => x"08782e81",
  1384 => x"b838778f",
  1385 => x"06a01757",
  1386 => x"54739138",
  1387 => x"80c6bc52",
  1388 => x"76518117",
  1389 => x"579eba2d",
  1390 => x"80c6bc56",
  1391 => x"807680f5",
  1392 => x"2d565474",
  1393 => x"742e8338",
  1394 => x"81547481",
  1395 => x"e52e80fd",
  1396 => x"38817075",
  1397 => x"06555c73",
  1398 => x"802e80f1",
  1399 => x"388b1680",
  1400 => x"f52d9806",
  1401 => x"597880e5",
  1402 => x"388b537c",
  1403 => x"5275519f",
  1404 => x"dd2d80c5",
  1405 => x"d40880d5",
  1406 => x"389c1608",
  1407 => x"51adf82d",
  1408 => x"80c5d408",
  1409 => x"841b0c9a",
  1410 => x"1680e02d",
  1411 => x"51aea92d",
  1412 => x"80c5d408",
  1413 => x"80c5d408",
  1414 => x"881c0c80",
  1415 => x"c5d40855",
  1416 => x"5580ccc8",
  1417 => x"08802e99",
  1418 => x"38941680",
  1419 => x"e02d51ae",
  1420 => x"a92d80c5",
  1421 => x"d408902b",
  1422 => x"83fff00a",
  1423 => x"06701651",
  1424 => x"5473881b",
  1425 => x"0c787a0c",
  1426 => x"7b54ad95",
  1427 => x"04811858",
  1428 => x"80cccc08",
  1429 => x"7826feca",
  1430 => x"3880ccc8",
  1431 => x"08802eb3",
  1432 => x"387a51a7",
  1433 => x"ce2d80c5",
  1434 => x"d40880c5",
  1435 => x"d40880ff",
  1436 => x"fffff806",
  1437 => x"555b7380",
  1438 => x"fffffff8",
  1439 => x"2e953880",
  1440 => x"c5d408fe",
  1441 => x"0580ccc0",
  1442 => x"082980cc",
  1443 => x"d4080557",
  1444 => x"ab970480",
  1445 => x"547380c5",
  1446 => x"d40c02b4",
  1447 => x"050d0402",
  1448 => x"f4050d74",
  1449 => x"70088105",
  1450 => x"710c7008",
  1451 => x"80ccc408",
  1452 => x"06535371",
  1453 => x"8f388813",
  1454 => x"0851a7ce",
  1455 => x"2d80c5d4",
  1456 => x"0888140c",
  1457 => x"810b80c5",
  1458 => x"d40c028c",
  1459 => x"050d0402",
  1460 => x"f0050d75",
  1461 => x"881108fe",
  1462 => x"0580ccc0",
  1463 => x"082980cc",
  1464 => x"d4081172",
  1465 => x"0880ccc4",
  1466 => x"08060579",
  1467 => x"55535454",
  1468 => x"9eba2d02",
  1469 => x"90050d04",
  1470 => x"02f4050d",
  1471 => x"7470882a",
  1472 => x"83fe8006",
  1473 => x"7072982a",
  1474 => x"0772882b",
  1475 => x"87fc8080",
  1476 => x"0673982b",
  1477 => x"81f00a06",
  1478 => x"71730707",
  1479 => x"80c5d40c",
  1480 => x"56515351",
  1481 => x"028c050d",
  1482 => x"0402f805",
  1483 => x"0d028e05",
  1484 => x"80f52d74",
  1485 => x"882b0770",
  1486 => x"83ffff06",
  1487 => x"80c5d40c",
  1488 => x"51028805",
  1489 => x"0d0402f4",
  1490 => x"050d7476",
  1491 => x"78535452",
  1492 => x"80712597",
  1493 => x"38727081",
  1494 => x"055480f5",
  1495 => x"2d727081",
  1496 => x"055481b7",
  1497 => x"2dff1151",
  1498 => x"70eb3880",
  1499 => x"7281b72d",
  1500 => x"028c050d",
  1501 => x"0402e805",
  1502 => x"0d775680",
  1503 => x"70565473",
  1504 => x"7624b638",
  1505 => x"80cccc08",
  1506 => x"742eae38",
  1507 => x"7351a8c7",
  1508 => x"2d80c5d4",
  1509 => x"0880c5d4",
  1510 => x"08098105",
  1511 => x"7080c5d4",
  1512 => x"08079f2a",
  1513 => x"77058117",
  1514 => x"57575353",
  1515 => x"74762489",
  1516 => x"3880cccc",
  1517 => x"087426d4",
  1518 => x"387280c5",
  1519 => x"d40c0298",
  1520 => x"050d0402",
  1521 => x"f0050d80",
  1522 => x"c5d00816",
  1523 => x"51aef52d",
  1524 => x"80c5d408",
  1525 => x"802e9f38",
  1526 => x"8b5380c5",
  1527 => x"d4085280",
  1528 => x"cabc51ae",
  1529 => x"c62d80cc",
  1530 => x"f8085473",
  1531 => x"802e8738",
  1532 => x"80cabc51",
  1533 => x"732d0290",
  1534 => x"050d0402",
  1535 => x"dc050d80",
  1536 => x"705a5574",
  1537 => x"80c5d008",
  1538 => x"25b43880",
  1539 => x"cccc0875",
  1540 => x"2eac3878",
  1541 => x"51a8c72d",
  1542 => x"80c5d408",
  1543 => x"09810570",
  1544 => x"80c5d408",
  1545 => x"079f2a76",
  1546 => x"05811b5b",
  1547 => x"56547480",
  1548 => x"c5d00825",
  1549 => x"893880cc",
  1550 => x"cc087926",
  1551 => x"d6388055",
  1552 => x"7880cccc",
  1553 => x"082781db",
  1554 => x"387851a8",
  1555 => x"c72d80c5",
  1556 => x"d408802e",
  1557 => x"81ad3880",
  1558 => x"c5d4088b",
  1559 => x"0580f52d",
  1560 => x"70842a70",
  1561 => x"81067710",
  1562 => x"78842b80",
  1563 => x"cabc0b80",
  1564 => x"f52d5c5c",
  1565 => x"53515556",
  1566 => x"73802e80",
  1567 => x"cb387416",
  1568 => x"822bb2c7",
  1569 => x"0b80c4a4",
  1570 => x"120c5477",
  1571 => x"75311080",
  1572 => x"ccfc1155",
  1573 => x"56907470",
  1574 => x"81055681",
  1575 => x"b72da074",
  1576 => x"81b72d76",
  1577 => x"81ff0681",
  1578 => x"16585473",
  1579 => x"802e8a38",
  1580 => x"9c5380ca",
  1581 => x"bc52b1c0",
  1582 => x"048b5380",
  1583 => x"c5d40852",
  1584 => x"80ccfe16",
  1585 => x"51b1fb04",
  1586 => x"7416822b",
  1587 => x"afc30b80",
  1588 => x"c4a4120c",
  1589 => x"547681ff",
  1590 => x"06811658",
  1591 => x"5473802e",
  1592 => x"8a389c53",
  1593 => x"80cabc52",
  1594 => x"b1f2048b",
  1595 => x"5380c5d4",
  1596 => x"08527775",
  1597 => x"311080cc",
  1598 => x"fc055176",
  1599 => x"55aec62d",
  1600 => x"b2980474",
  1601 => x"90297531",
  1602 => x"701080cc",
  1603 => x"fc055154",
  1604 => x"80c5d408",
  1605 => x"7481b72d",
  1606 => x"81195974",
  1607 => x"8b24a338",
  1608 => x"b0c00474",
  1609 => x"90297531",
  1610 => x"701080cc",
  1611 => x"fc058c77",
  1612 => x"31575154",
  1613 => x"807481b7",
  1614 => x"2d9e14ff",
  1615 => x"16565474",
  1616 => x"f33802a4",
  1617 => x"050d0402",
  1618 => x"fc050d80",
  1619 => x"c5d00813",
  1620 => x"51aef52d",
  1621 => x"80c5d408",
  1622 => x"802e8938",
  1623 => x"80c5d408",
  1624 => x"51a09c2d",
  1625 => x"800b80c5",
  1626 => x"d00caffb",
  1627 => x"2d91832d",
  1628 => x"0284050d",
  1629 => x"0402fc05",
  1630 => x"0d725170",
  1631 => x"fd2eb038",
  1632 => x"70fd248a",
  1633 => x"3870fc2e",
  1634 => x"80cc38b3",
  1635 => x"e00470fe",
  1636 => x"2eb73870",
  1637 => x"ff2e0981",
  1638 => x"0680c538",
  1639 => x"80c5d008",
  1640 => x"5170802e",
  1641 => x"bb38ff11",
  1642 => x"80c5d00c",
  1643 => x"b3e00480",
  1644 => x"c5d008f0",
  1645 => x"057080c5",
  1646 => x"d00c5170",
  1647 => x"8025a138",
  1648 => x"800b80c5",
  1649 => x"d00cb3e0",
  1650 => x"0480c5d0",
  1651 => x"08810580",
  1652 => x"c5d00cb3",
  1653 => x"e00480c5",
  1654 => x"d0089005",
  1655 => x"80c5d00c",
  1656 => x"affb2d91",
  1657 => x"832d0284",
  1658 => x"050d0402",
  1659 => x"fc050d80",
  1660 => x"0b80c5d0",
  1661 => x"0caffb2d",
  1662 => x"90932d80",
  1663 => x"c5d40880",
  1664 => x"c5c00c80",
  1665 => x"c49c5192",
  1666 => x"a62d0284",
  1667 => x"050d0471",
  1668 => x"80ccf80c",
  1669 => x"04000000",
  1670 => x"00ffffff",
  1671 => x"ff00ffff",
  1672 => x"ffff00ff",
  1673 => x"ffffff00",
  1674 => x"45786974",
  1675 => x"00000000",
  1676 => x"506f7420",
  1677 => x"33263420",
  1678 => x"4a6f7920",
  1679 => x"32204669",
  1680 => x"72652032",
  1681 => x"2f330000",
  1682 => x"506f7420",
  1683 => x"33263420",
  1684 => x"4d6f7573",
  1685 => x"65000000",
  1686 => x"506f7420",
  1687 => x"33263420",
  1688 => x"50616464",
  1689 => x"6c657320",
  1690 => x"33263400",
  1691 => x"506f7420",
  1692 => x"31263220",
  1693 => x"4a6f7920",
  1694 => x"31204669",
  1695 => x"72652032",
  1696 => x"2f330000",
  1697 => x"506f7420",
  1698 => x"31263220",
  1699 => x"4d6f7573",
  1700 => x"65000000",
  1701 => x"506f7420",
  1702 => x"31263220",
  1703 => x"50616464",
  1704 => x"6c657320",
  1705 => x"31263200",
  1706 => x"506f7274",
  1707 => x"20554152",
  1708 => x"54000000",
  1709 => x"506f7274",
  1710 => x"204a6f79",
  1711 => x"73746963",
  1712 => x"6b730000",
  1713 => x"4a6f7973",
  1714 => x"7469636b",
  1715 => x"73204e6f",
  1716 => x"726d616c",
  1717 => x"00000000",
  1718 => x"4a6f7973",
  1719 => x"7469636b",
  1720 => x"73207377",
  1721 => x"61707065",
  1722 => x"64000000",
  1723 => x"44696769",
  1724 => x"6d617820",
  1725 => x"4e6f0000",
  1726 => x"44696769",
  1727 => x"6d617820",
  1728 => x"24444530",
  1729 => x"30000000",
  1730 => x"44696769",
  1731 => x"6d617820",
  1732 => x"24444630",
  1733 => x"30000000",
  1734 => x"53746572",
  1735 => x"656f206d",
  1736 => x"6978204e",
  1737 => x"6f000000",
  1738 => x"53746572",
  1739 => x"656f206d",
  1740 => x"69782032",
  1741 => x"35250000",
  1742 => x"53746572",
  1743 => x"656f206d",
  1744 => x"69782035",
  1745 => x"30250000",
  1746 => x"53746572",
  1747 => x"656f206d",
  1748 => x"69782031",
  1749 => x"30302500",
  1750 => x"536f756e",
  1751 => x"64206578",
  1752 => x"70616e73",
  1753 => x"696f6e20",
  1754 => x"4e6f0000",
  1755 => x"536f756e",
  1756 => x"64206578",
  1757 => x"70616e73",
  1758 => x"696f6e20",
  1759 => x"4f504c32",
  1760 => x"00000000",
  1761 => x"53494420",
  1762 => x"72696768",
  1763 => x"74204164",
  1764 => x"64722053",
  1765 => x"616d6500",
  1766 => x"53494420",
  1767 => x"72696768",
  1768 => x"74204164",
  1769 => x"64722024",
  1770 => x"44343230",
  1771 => x"00000000",
  1772 => x"53494420",
  1773 => x"72696768",
  1774 => x"74204164",
  1775 => x"64722024",
  1776 => x"44353030",
  1777 => x"00000000",
  1778 => x"53494420",
  1779 => x"52696768",
  1780 => x"74203635",
  1781 => x"38310000",
  1782 => x"53494420",
  1783 => x"52696768",
  1784 => x"74203835",
  1785 => x"38300000",
  1786 => x"53494420",
  1787 => x"4c656674",
  1788 => x"20363538",
  1789 => x"31000000",
  1790 => x"53494420",
  1791 => x"4c656674",
  1792 => x"20383538",
  1793 => x"30000000",
  1794 => x"50616c65",
  1795 => x"74746520",
  1796 => x"43363400",
  1797 => x"50616c65",
  1798 => x"74746520",
  1799 => x"43655065",
  1800 => x"43655261",
  1801 => x"00000000",
  1802 => x"50616c65",
  1803 => x"74746520",
  1804 => x"50657074",
  1805 => x"6f000000",
  1806 => x"50616c65",
  1807 => x"74746520",
  1808 => x"436f6d75",
  1809 => x"6e697479",
  1810 => x"00000000",
  1811 => x"5363616e",
  1812 => x"646f7562",
  1813 => x"6c657220",
  1814 => x"4e6f6e65",
  1815 => x"00000000",
  1816 => x"5363616e",
  1817 => x"646f7562",
  1818 => x"6c657220",
  1819 => x"43525420",
  1820 => x"32352500",
  1821 => x"5363616e",
  1822 => x"646f7562",
  1823 => x"6c657220",
  1824 => x"43525420",
  1825 => x"35302500",
  1826 => x"5363616e",
  1827 => x"646f7562",
  1828 => x"6c657220",
  1829 => x"43525420",
  1830 => x"37352500",
  1831 => x"4f726967",
  1832 => x"696e616c",
  1833 => x"20666f72",
  1834 => x"6d617400",
  1835 => x"46756c6c",
  1836 => x"20736372",
  1837 => x"65656e00",
  1838 => x"466f726d",
  1839 => x"6174205b",
  1840 => x"41524331",
  1841 => x"5d000000",
  1842 => x"466f726d",
  1843 => x"6174205b",
  1844 => x"41524332",
  1845 => x"5d000000",
  1846 => x"4f726967",
  1847 => x"696e616c",
  1848 => x"20617370",
  1849 => x"65637420",
  1850 => x"72617469",
  1851 => x"6f000000",
  1852 => x"57696465",
  1853 => x"20617370",
  1854 => x"65637420",
  1855 => x"72617469",
  1856 => x"6f000000",
  1857 => x"56696465",
  1858 => x"6f205041",
  1859 => x"4c000000",
  1860 => x"56696465",
  1861 => x"6f204e54",
  1862 => x"53430000",
  1863 => x"2020203d",
  1864 => x"20434f4d",
  1865 => x"4f444f52",
  1866 => x"45202036",
  1867 => x"34203d20",
  1868 => x"20200000",
  1869 => x"20202020",
  1870 => x"20204e65",
  1871 => x"75726f52",
  1872 => x"756c657a",
  1873 => x"20202020",
  1874 => x"20200000",
  1875 => x"20202020",
  1876 => x"20202020",
  1877 => x"20202020",
  1878 => x"20202020",
  1879 => x"20202020",
  1880 => x"20200000",
  1881 => x"52657365",
  1882 => x"74000000",
  1883 => x"52657365",
  1884 => x"74202620",
  1885 => x"44657461",
  1886 => x"63682063",
  1887 => x"61727472",
  1888 => x"69646765",
  1889 => x"00000000",
  1890 => x"56696465",
  1891 => x"6f201000",
  1892 => x"41756469",
  1893 => x"6f201000",
  1894 => x"50756572",
  1895 => x"746f7320",
  1896 => x"10000000",
  1897 => x"456a6563",
  1898 => x"74207461",
  1899 => x"70650000",
  1900 => x"506c6179",
  1901 => x"2f53746f",
  1902 => x"70205461",
  1903 => x"70650000",
  1904 => x"4c6f6164",
  1905 => x"20446973",
  1906 => x"6b2f5461",
  1907 => x"70652f43",
  1908 => x"61727420",
  1909 => x"10000000",
  1910 => x"4469736b",
  1911 => x"20777269",
  1912 => x"7465204f",
  1913 => x"6e000000",
  1914 => x"4469736b",
  1915 => x"20777269",
  1916 => x"7465204f",
  1917 => x"66660000",
  1918 => x"54617065",
  1919 => x"20736f75",
  1920 => x"6e64204f",
  1921 => x"66660000",
  1922 => x"54617065",
  1923 => x"20736f75",
  1924 => x"6e64204f",
  1925 => x"6e000000",
  1926 => x"4b65726e",
  1927 => x"656c206c",
  1928 => x"6f616461",
  1929 => x"626c6500",
  1930 => x"4b65726e",
  1931 => x"656c2043",
  1932 => x"36340000",
  1933 => x"4b65726e",
  1934 => x"656c2043",
  1935 => x"36344753",
  1936 => x"00000000",
  1937 => x"4b65726e",
  1938 => x"656c204a",
  1939 => x"6170616e",
  1940 => x"00000000",
  1941 => x"43617267",
  1942 => x"61204661",
  1943 => x"6c6c6964",
  1944 => x"61000000",
  1945 => x"4f4b0000",
  1946 => x"16200000",
  1947 => x"14200000",
  1948 => x"15200000",
  1949 => x"53442069",
  1950 => x"6e69742e",
  1951 => x"2e2e0a00",
  1952 => x"53442063",
  1953 => x"61726420",
  1954 => x"72657365",
  1955 => x"74206661",
  1956 => x"696c6564",
  1957 => x"210a0000",
  1958 => x"53444843",
  1959 => x"20657272",
  1960 => x"6f72210a",
  1961 => x"00000000",
  1962 => x"57726974",
  1963 => x"65206661",
  1964 => x"696c6564",
  1965 => x"0a000000",
  1966 => x"52656164",
  1967 => x"20666169",
  1968 => x"6c65640a",
  1969 => x"00000000",
  1970 => x"43617264",
  1971 => x"20696e69",
  1972 => x"74206661",
  1973 => x"696c6564",
  1974 => x"0a000000",
  1975 => x"46415431",
  1976 => x"36202020",
  1977 => x"00000000",
  1978 => x"46415433",
  1979 => x"32202020",
  1980 => x"00000000",
  1981 => x"4e6f2070",
  1982 => x"61727469",
  1983 => x"74696f6e",
  1984 => x"20736967",
  1985 => x"0a000000",
  1986 => x"42616420",
  1987 => x"70617274",
  1988 => x"0a000000",
  1989 => x"4261636b",
  1990 => x"00000000",
  1991 => x"00000002",
  1992 => x"00000003",
  1993 => x"00001f88",
  1994 => x"00000002",
  1995 => x"00000003",
  1996 => x"00001f80",
  1997 => x"00000002",
  1998 => x"00000003",
  1999 => x"00001f74",
  2000 => x"00000003",
  2001 => x"00000003",
  2002 => x"00001f68",
  2003 => x"00000003",
  2004 => x"00000004",
  2005 => x"00001a28",
  2006 => x"000020c4",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00000000",
  2010 => x"00001a30",
  2011 => x"00001a48",
  2012 => x"00001a58",
  2013 => x"00001a6c",
  2014 => x"00001a84",
  2015 => x"00001a94",
  2016 => x"00001aa8",
  2017 => x"00001ab4",
  2018 => x"00001ac4",
  2019 => x"00001ad8",
  2020 => x"00000003",
  2021 => x"00002028",
  2022 => x"00000002",
  2023 => x"00000003",
  2024 => x"00002020",
  2025 => x"00000002",
  2026 => x"00000003",
  2027 => x"00002014",
  2028 => x"00000003",
  2029 => x"00000003",
  2030 => x"0000200c",
  2031 => x"00000002",
  2032 => x"00000003",
  2033 => x"00001ffc",
  2034 => x"00000004",
  2035 => x"00000003",
  2036 => x"00001ff0",
  2037 => x"00000003",
  2038 => x"00000004",
  2039 => x"00001a28",
  2040 => x"000020c4",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00001aec",
  2045 => x"00001af8",
  2046 => x"00001b08",
  2047 => x"00001b18",
  2048 => x"00001b28",
  2049 => x"00001b38",
  2050 => x"00001b48",
  2051 => x"00001b58",
  2052 => x"00001b6c",
  2053 => x"00001b84",
  2054 => x"00001b98",
  2055 => x"00001bb0",
  2056 => x"00001bc8",
  2057 => x"00001bd8",
  2058 => x"00001be8",
  2059 => x"00001bf8",
  2060 => x"00000003",
  2061 => x"000020bc",
  2062 => x"00000002",
  2063 => x"00000003",
  2064 => x"000020b4",
  2065 => x"00000002",
  2066 => x"00000003",
  2067 => x"000020a4",
  2068 => x"00000004",
  2069 => x"00000003",
  2070 => x"00002094",
  2071 => x"00000004",
  2072 => x"00000003",
  2073 => x"00002084",
  2074 => x"00000004",
  2075 => x"00000004",
  2076 => x"00001a28",
  2077 => x"000020c4",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00001c08",
  2082 => x"00001c14",
  2083 => x"00001c28",
  2084 => x"00001c38",
  2085 => x"00001c4c",
  2086 => x"00001c60",
  2087 => x"00001c74",
  2088 => x"00001c88",
  2089 => x"00001c9c",
  2090 => x"00001cac",
  2091 => x"00001cb8",
  2092 => x"00001cc8",
  2093 => x"00001cd8",
  2094 => x"00001cf0",
  2095 => x"00001d04",
  2096 => x"00001d10",
  2097 => x"00000002",
  2098 => x"00001d1c",
  2099 => x"00000000",
  2100 => x"00000002",
  2101 => x"00001d34",
  2102 => x"00000000",
  2103 => x"00000002",
  2104 => x"00001d4c",
  2105 => x"00000000",
  2106 => x"00000002",
  2107 => x"00001d64",
  2108 => x"00000371",
  2109 => x"00000002",
  2110 => x"00001d6c",
  2111 => x"00000388",
  2112 => x"00000004",
  2113 => x"00001d88",
  2114 => x"00002030",
  2115 => x"00000004",
  2116 => x"00001d90",
  2117 => x"00001f90",
  2118 => x"00000004",
  2119 => x"00001d98",
  2120 => x"00001f20",
  2121 => x"00000003",
  2122 => x"00002194",
  2123 => x"00000004",
  2124 => x"00000003",
  2125 => x"0000218c",
  2126 => x"00000002",
  2127 => x"00000003",
  2128 => x"00002184",
  2129 => x"00000002",
  2130 => x"00000002",
  2131 => x"00001da4",
  2132 => x"000003b8",
  2133 => x"00000002",
  2134 => x"00001db0",
  2135 => x"000003a0",
  2136 => x"00000002",
  2137 => x"00001dc0",
  2138 => x"000019eb",
  2139 => x"00000002",
  2140 => x"00001a28",
  2141 => x"0000081c",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00001dd8",
  2146 => x"00001de8",
  2147 => x"00001df8",
  2148 => x"00001e08",
  2149 => x"00001e18",
  2150 => x"00001e28",
  2151 => x"00001e34",
  2152 => x"00001e44",
  2153 => x"00000004",
  2154 => x"00001e54",
  2155 => x"000021a4",
  2156 => x"00000004",
  2157 => x"00001e64",
  2158 => x"000020c4",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000002",
  2184 => x"0000267c",
  2185 => x"000017c3",
  2186 => x"00000002",
  2187 => x"0000269a",
  2188 => x"000017c3",
  2189 => x"00000002",
  2190 => x"000026b8",
  2191 => x"000017c3",
  2192 => x"00000002",
  2193 => x"000026d6",
  2194 => x"000017c3",
  2195 => x"00000002",
  2196 => x"000026f4",
  2197 => x"000017c3",
  2198 => x"00000002",
  2199 => x"00002712",
  2200 => x"000017c3",
  2201 => x"00000002",
  2202 => x"00002730",
  2203 => x"000017c3",
  2204 => x"00000002",
  2205 => x"0000274e",
  2206 => x"000017c3",
  2207 => x"00000002",
  2208 => x"0000276c",
  2209 => x"000017c3",
  2210 => x"00000002",
  2211 => x"0000278a",
  2212 => x"000017c3",
  2213 => x"00000002",
  2214 => x"000027a8",
  2215 => x"000017c3",
  2216 => x"00000002",
  2217 => x"000027c6",
  2218 => x"000017c3",
  2219 => x"00000002",
  2220 => x"000027e4",
  2221 => x"000017c3",
  2222 => x"00000004",
  2223 => x"00001f14",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00001975",
  2228 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

