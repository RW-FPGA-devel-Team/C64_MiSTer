-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c6",
     9 => x"b4080b0b",
    10 => x"80c6b808",
    11 => x"0b0b80c6",
    12 => x"bc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c6bc0c0b",
    16 => x"0b80c6b8",
    17 => x"0c0b0b80",
    18 => x"c6b40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb4ac",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c6b470",
    57 => x"80d0e427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5189dd",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c6",
    65 => x"c40c9f0b",
    66 => x"80c6c80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c6c808ff",
    70 => x"0580c6c8",
    71 => x"0c80c6c8",
    72 => x"088025e8",
    73 => x"3880c6c4",
    74 => x"08ff0580",
    75 => x"c6c40c80",
    76 => x"c6c40880",
    77 => x"25d03880",
    78 => x"0b80c6c8",
    79 => x"0c800b80",
    80 => x"c6c40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c6c408",
   100 => x"25913882",
   101 => x"c82d80c6",
   102 => x"c408ff05",
   103 => x"80c6c40c",
   104 => x"838a0480",
   105 => x"c6c40880",
   106 => x"c6c80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c6c408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c6c80881",
   116 => x"0580c6c8",
   117 => x"0c80c6c8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c6c8",
   121 => x"0c80c6c4",
   122 => x"08810580",
   123 => x"c6c40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c6",
   128 => x"c8088105",
   129 => x"80c6c80c",
   130 => x"80c6c808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c6c8",
   134 => x"0c80c6c4",
   135 => x"08810580",
   136 => x"c6c40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"c6cc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"c6cc0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280c6",
   177 => x"cc088407",
   178 => x"80c6cc0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b0bbe",
   183 => x"fc0c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80c6cc",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80c6",
   208 => x"b40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050d84bf",
   216 => x"5186c72d",
   217 => x"ff115170",
   218 => x"8025f638",
   219 => x"0284050d",
   220 => x"0402fc05",
   221 => x"0dec5183",
   222 => x"710c86c7",
   223 => x"2d82710c",
   224 => x"90b12d02",
   225 => x"84050d04",
   226 => x"02fc050d",
   227 => x"ec518182",
   228 => x"710c86c7",
   229 => x"2d82710c",
   230 => x"90b12d02",
   231 => x"84050d04",
   232 => x"02fc050d",
   233 => x"ec5180c2",
   234 => x"710c86c7",
   235 => x"2d82710c",
   236 => x"90b12d02",
   237 => x"84050d04",
   238 => x"02fc050d",
   239 => x"ec518282",
   240 => x"710c86c7",
   241 => x"2d82710c",
   242 => x"90b12d02",
   243 => x"84050d04",
   244 => x"02fc050d",
   245 => x"ec519271",
   246 => x"0c86c72d",
   247 => x"82710c02",
   248 => x"84050d04",
   249 => x"02d0050d",
   250 => x"7d548074",
   251 => x"5380c6d0",
   252 => x"525bab97",
   253 => x"2d80c6b4",
   254 => x"087b2e81",
   255 => x"b63880c6",
   256 => x"d40870f8",
   257 => x"0c891580",
   258 => x"f52d8a16",
   259 => x"80f52d71",
   260 => x"82802905",
   261 => x"881780f5",
   262 => x"2d708480",
   263 => x"802912f4",
   264 => x"0c575556",
   265 => x"58a40bec",
   266 => x"0c7aff19",
   267 => x"585a767b",
   268 => x"2e8b3881",
   269 => x"1a77812a",
   270 => x"585a76f7",
   271 => x"38f71a5a",
   272 => x"815b8078",
   273 => x"2580ec38",
   274 => x"79527651",
   275 => x"84a82d80",
   276 => x"c79c5280",
   277 => x"c6d051ad",
   278 => x"e42d80c6",
   279 => x"b408802e",
   280 => x"b93880c7",
   281 => x"9c5c83fc",
   282 => x"597b7084",
   283 => x"055d0870",
   284 => x"81ff0671",
   285 => x"882a7081",
   286 => x"ff067390",
   287 => x"2a7081ff",
   288 => x"0675982a",
   289 => x"e80ce80c",
   290 => x"58e80c57",
   291 => x"e80cfc1a",
   292 => x"5a537880",
   293 => x"25d33889",
   294 => x"a20480c6",
   295 => x"b4085b84",
   296 => x"805880c6",
   297 => x"d051adb4",
   298 => x"2dfc8018",
   299 => x"81185858",
   300 => x"88c20486",
   301 => x"da2d840b",
   302 => x"ec0c7a80",
   303 => x"2e8e3880",
   304 => x"c2a45192",
   305 => x"bb2d90b1",
   306 => x"2d89d304",
   307 => x"80c48451",
   308 => x"92bb2d7a",
   309 => x"80c6b40c",
   310 => x"02b0050d",
   311 => x"0402ec05",
   312 => x"0d840bec",
   313 => x"0c908f2d",
   314 => x"8ce12d81",
   315 => x"f92da1d7",
   316 => x"2d80c6b4",
   317 => x"08802e82",
   318 => x"d13887e4",
   319 => x"51b4a42d",
   320 => x"80c2a451",
   321 => x"92bb2d90",
   322 => x"b12d8ced",
   323 => x"2d92ce2d",
   324 => x"80c1980b",
   325 => x"80f52d70",
   326 => x"822b8406",
   327 => x"80c1a40b",
   328 => x"80f52d70",
   329 => x"982b8180",
   330 => x"0a0680c1",
   331 => x"b00b80f5",
   332 => x"2d70842b",
   333 => x"b0067473",
   334 => x"070780c1",
   335 => x"bc0b80f5",
   336 => x"2d70882b",
   337 => x"86800680",
   338 => x"c1c80b80",
   339 => x"f52d7372",
   340 => x"07719e2b",
   341 => x"07bff80b",
   342 => x"80f52d70",
   343 => x"8d2b80c0",
   344 => x"800680c0",
   345 => x"840b80f5",
   346 => x"2d70902b",
   347 => x"84808006",
   348 => x"74730707",
   349 => x"80c0900b",
   350 => x"80f52d70",
   351 => x"962b8680",
   352 => x"0a0680c0",
   353 => x"9c0b80f5",
   354 => x"2d708c2b",
   355 => x"a0800674",
   356 => x"73070780",
   357 => x"c0a80b80",
   358 => x"f52d7092",
   359 => x"2bb08080",
   360 => x"0680c0b4",
   361 => x"0b80f52d",
   362 => x"70942b98",
   363 => x"800a0674",
   364 => x"730707bf",
   365 => x"880b80f5",
   366 => x"2d70832b",
   367 => x"8806bf94",
   368 => x"0b80f52d",
   369 => x"70108206",
   370 => x"74730707",
   371 => x"bfa00b80",
   372 => x"f52d709a",
   373 => x"2bb00a06",
   374 => x"bfac0b80",
   375 => x"f52d709c",
   376 => x"2b8c0a06",
   377 => x"74730707",
   378 => x"80c38c0b",
   379 => x"80f52d70",
   380 => x"8e2b8380",
   381 => x"800680c3",
   382 => x"980b80f5",
   383 => x"2d708b2b",
   384 => x"90800674",
   385 => x"73070780",
   386 => x"c3a40b80",
   387 => x"f52d7081",
   388 => x"06a02b72",
   389 => x"07fc0c53",
   390 => x"54545454",
   391 => x"54545454",
   392 => x"54545454",
   393 => x"54545454",
   394 => x"54545454",
   395 => x"54545553",
   396 => x"54545753",
   397 => x"54525757",
   398 => x"53538652",
   399 => x"80c6b408",
   400 => x"83388452",
   401 => x"71ec0c8a",
   402 => x"8a04800b",
   403 => x"80c6b40c",
   404 => x"0294050d",
   405 => x"0471980c",
   406 => x"04ffb008",
   407 => x"80c6b40c",
   408 => x"04810bff",
   409 => x"b00c0480",
   410 => x"0bffb00c",
   411 => x"0402f405",
   412 => x"0d8dfb04",
   413 => x"80c6b408",
   414 => x"81f02e09",
   415 => x"81068a38",
   416 => x"810b80c4",
   417 => x"e80c8dfb",
   418 => x"0480c6b4",
   419 => x"0881e02e",
   420 => x"0981068a",
   421 => x"38810b80",
   422 => x"c4ec0c8d",
   423 => x"fb0480c6",
   424 => x"b4085280",
   425 => x"c4ec0880",
   426 => x"2e893880",
   427 => x"c6b40881",
   428 => x"80055271",
   429 => x"842c728f",
   430 => x"06535380",
   431 => x"c4e80880",
   432 => x"2e9a3872",
   433 => x"842980c4",
   434 => x"a8057213",
   435 => x"81712b70",
   436 => x"09730806",
   437 => x"730c5153",
   438 => x"538def04",
   439 => x"72842980",
   440 => x"c4a80572",
   441 => x"1383712b",
   442 => x"72080772",
   443 => x"0c535380",
   444 => x"0b80c4ec",
   445 => x"0c800b80",
   446 => x"c4e80c80",
   447 => x"c6dc518f",
   448 => x"822d80c6",
   449 => x"b408ff24",
   450 => x"feea3880",
   451 => x"0b80c6b4",
   452 => x"0c028c05",
   453 => x"0d0402f8",
   454 => x"050d80c4",
   455 => x"a8528f51",
   456 => x"80727084",
   457 => x"05540cff",
   458 => x"11517080",
   459 => x"25f23802",
   460 => x"88050d04",
   461 => x"02f0050d",
   462 => x"75518ce7",
   463 => x"2d70822c",
   464 => x"fc0680c4",
   465 => x"a8117210",
   466 => x"9e067108",
   467 => x"70722a70",
   468 => x"83068274",
   469 => x"2b700974",
   470 => x"06760c54",
   471 => x"51565753",
   472 => x"51538ce1",
   473 => x"2d7180c6",
   474 => x"b40c0290",
   475 => x"050d0402",
   476 => x"fc050d72",
   477 => x"5180710c",
   478 => x"800b8412",
   479 => x"0c028405",
   480 => x"0d0402f0",
   481 => x"050d7570",
   482 => x"08841208",
   483 => x"535353ff",
   484 => x"5471712e",
   485 => x"a8388ce7",
   486 => x"2d841308",
   487 => x"70842914",
   488 => x"88117008",
   489 => x"7081ff06",
   490 => x"84180881",
   491 => x"11870684",
   492 => x"1a0c5351",
   493 => x"55515151",
   494 => x"8ce12d71",
   495 => x"547380c6",
   496 => x"b40c0290",
   497 => x"050d0402",
   498 => x"f8050d8c",
   499 => x"e72de008",
   500 => x"708b2a70",
   501 => x"81065152",
   502 => x"5270802e",
   503 => x"a13880c6",
   504 => x"dc087084",
   505 => x"2980c6e4",
   506 => x"057381ff",
   507 => x"06710c51",
   508 => x"5180c6dc",
   509 => x"08811187",
   510 => x"0680c6dc",
   511 => x"0c51800b",
   512 => x"80c7840c",
   513 => x"8cd92d8c",
   514 => x"e12d0288",
   515 => x"050d0402",
   516 => x"fc050d80",
   517 => x"c6dc518e",
   518 => x"ef2d8e96",
   519 => x"2d8fc751",
   520 => x"8cd52d02",
   521 => x"84050d04",
   522 => x"80c78808",
   523 => x"80c6b40c",
   524 => x"0402fc05",
   525 => x"0d90bb04",
   526 => x"8ced2d80",
   527 => x"f6518eb4",
   528 => x"2d80c6b4",
   529 => x"08f23880",
   530 => x"da518eb4",
   531 => x"2d80c6b4",
   532 => x"08e63880",
   533 => x"c6b40880",
   534 => x"c4f40c80",
   535 => x"c6b40851",
   536 => x"858d2d02",
   537 => x"84050d04",
   538 => x"02ec050d",
   539 => x"76548052",
   540 => x"870b8815",
   541 => x"80f52d56",
   542 => x"53747224",
   543 => x"8338a053",
   544 => x"72518384",
   545 => x"2d81128b",
   546 => x"1580f52d",
   547 => x"54527272",
   548 => x"25de3802",
   549 => x"94050d04",
   550 => x"02f0050d",
   551 => x"80c78808",
   552 => x"5481f92d",
   553 => x"800b80c7",
   554 => x"8c0c7308",
   555 => x"802e8186",
   556 => x"38820b80",
   557 => x"c6c80c80",
   558 => x"c78c088f",
   559 => x"0680c6c4",
   560 => x"0c730852",
   561 => x"71832e96",
   562 => x"38718326",
   563 => x"89387181",
   564 => x"2eaf3892",
   565 => x"9f047185",
   566 => x"2e9f3892",
   567 => x"9f048814",
   568 => x"80f52d84",
   569 => x"1508bdc8",
   570 => x"53545286",
   571 => x"a02d7184",
   572 => x"29137008",
   573 => x"525292a3",
   574 => x"04735190",
   575 => x"e82d929f",
   576 => x"0480c4f0",
   577 => x"08881508",
   578 => x"2c708106",
   579 => x"51527180",
   580 => x"2e8738bd",
   581 => x"cc51929c",
   582 => x"04bdd051",
   583 => x"86a02d84",
   584 => x"14085186",
   585 => x"a02d80c7",
   586 => x"8c088105",
   587 => x"80c78c0c",
   588 => x"8c145491",
   589 => x"aa040290",
   590 => x"050d0471",
   591 => x"80c7880c",
   592 => x"91982d80",
   593 => x"c78c08ff",
   594 => x"0580c790",
   595 => x"0c0402e8",
   596 => x"050d80c7",
   597 => x"880880c7",
   598 => x"94085755",
   599 => x"87518eb4",
   600 => x"2d80c6b4",
   601 => x"08812a70",
   602 => x"81065152",
   603 => x"71802ea3",
   604 => x"3892f704",
   605 => x"8ced2d87",
   606 => x"518eb42d",
   607 => x"80c6b408",
   608 => x"f33880c4",
   609 => x"f4088132",
   610 => x"7080c4f4",
   611 => x"0c705252",
   612 => x"858d2d80",
   613 => x"fe518eb4",
   614 => x"2d80c6b4",
   615 => x"08802ea9",
   616 => x"3880c4f4",
   617 => x"08802e92",
   618 => x"38800b80",
   619 => x"c4f40c80",
   620 => x"51858d2d",
   621 => x"93ba048c",
   622 => x"ed2d80fe",
   623 => x"518eb42d",
   624 => x"80c6b408",
   625 => x"f23887d0",
   626 => x"2d80c4f4",
   627 => x"08903881",
   628 => x"fd518eb4",
   629 => x"2d81fa51",
   630 => x"8eb42d99",
   631 => x"b30481f5",
   632 => x"518eb42d",
   633 => x"80c6b408",
   634 => x"812a7081",
   635 => x"06515271",
   636 => x"802eb338",
   637 => x"80c79008",
   638 => x"5271802e",
   639 => x"8a38ff12",
   640 => x"80c7900c",
   641 => x"94a60480",
   642 => x"c78c0810",
   643 => x"80c78c08",
   644 => x"05708429",
   645 => x"16515288",
   646 => x"1208802e",
   647 => x"8938ff51",
   648 => x"88120852",
   649 => x"712d81f2",
   650 => x"518eb42d",
   651 => x"80c6b408",
   652 => x"812a7081",
   653 => x"06515271",
   654 => x"802eb438",
   655 => x"80c78c08",
   656 => x"ff1180c7",
   657 => x"90085653",
   658 => x"53737225",
   659 => x"8a388114",
   660 => x"80c7900c",
   661 => x"94ef0472",
   662 => x"10137084",
   663 => x"29165152",
   664 => x"88120880",
   665 => x"2e8938fe",
   666 => x"51881208",
   667 => x"52712d81",
   668 => x"fd518eb4",
   669 => x"2d80c6b4",
   670 => x"08812a70",
   671 => x"81065152",
   672 => x"71802eb1",
   673 => x"3880c790",
   674 => x"08802e8a",
   675 => x"38800b80",
   676 => x"c7900c95",
   677 => x"b50480c7",
   678 => x"8c081080",
   679 => x"c78c0805",
   680 => x"70842916",
   681 => x"51528812",
   682 => x"08802e89",
   683 => x"38fd5188",
   684 => x"12085271",
   685 => x"2d81fa51",
   686 => x"8eb42d80",
   687 => x"c6b40881",
   688 => x"2a708106",
   689 => x"51527180",
   690 => x"2eb13880",
   691 => x"c78c08ff",
   692 => x"11545280",
   693 => x"c7900873",
   694 => x"25893872",
   695 => x"80c7900c",
   696 => x"95fb0471",
   697 => x"10127084",
   698 => x"29165152",
   699 => x"88120880",
   700 => x"2e8938fc",
   701 => x"51881208",
   702 => x"52712d80",
   703 => x"c7900870",
   704 => x"53547380",
   705 => x"2e8a388c",
   706 => x"15ff1555",
   707 => x"55968204",
   708 => x"820b80c6",
   709 => x"c80c718f",
   710 => x"0680c6c4",
   711 => x"0c81eb51",
   712 => x"8eb42d80",
   713 => x"c6b40881",
   714 => x"2a708106",
   715 => x"51527180",
   716 => x"2ead3874",
   717 => x"08852e09",
   718 => x"8106a438",
   719 => x"881580f5",
   720 => x"2dff0552",
   721 => x"71881681",
   722 => x"b72d7198",
   723 => x"2b527180",
   724 => x"25883880",
   725 => x"0b881681",
   726 => x"b72d7451",
   727 => x"90e82d81",
   728 => x"f4518eb4",
   729 => x"2d80c6b4",
   730 => x"08812a70",
   731 => x"81065152",
   732 => x"71802eb3",
   733 => x"38740885",
   734 => x"2e098106",
   735 => x"aa388815",
   736 => x"80f52d81",
   737 => x"05527188",
   738 => x"1681b72d",
   739 => x"7181ff06",
   740 => x"8b1680f5",
   741 => x"2d545272",
   742 => x"72278738",
   743 => x"72881681",
   744 => x"b72d7451",
   745 => x"90e82d80",
   746 => x"da518eb4",
   747 => x"2d80c6b4",
   748 => x"08812a70",
   749 => x"81065152",
   750 => x"71802e81",
   751 => x"ad3880c7",
   752 => x"880880c7",
   753 => x"90085553",
   754 => x"73802e8a",
   755 => x"388c13ff",
   756 => x"15555397",
   757 => x"c8047208",
   758 => x"5271822e",
   759 => x"a6387182",
   760 => x"26893871",
   761 => x"812eaa38",
   762 => x"98ea0471",
   763 => x"832eb438",
   764 => x"71842e09",
   765 => x"810680f2",
   766 => x"38881308",
   767 => x"5192bb2d",
   768 => x"98ea0480",
   769 => x"c7900851",
   770 => x"88130852",
   771 => x"712d98ea",
   772 => x"04810b88",
   773 => x"14082b80",
   774 => x"c4f00832",
   775 => x"80c4f00c",
   776 => x"98be0488",
   777 => x"1380f52d",
   778 => x"81058b14",
   779 => x"80f52d53",
   780 => x"54717424",
   781 => x"83388054",
   782 => x"73881481",
   783 => x"b72d9198",
   784 => x"2d98ea04",
   785 => x"7508802e",
   786 => x"a4387508",
   787 => x"518eb42d",
   788 => x"80c6b408",
   789 => x"81065271",
   790 => x"802e8c38",
   791 => x"80c79008",
   792 => x"51841608",
   793 => x"52712d88",
   794 => x"165675d8",
   795 => x"38805480",
   796 => x"0b80c6c8",
   797 => x"0c738f06",
   798 => x"80c6c40c",
   799 => x"a0527380",
   800 => x"c790082e",
   801 => x"09810699",
   802 => x"3880c78c",
   803 => x"08ff0574",
   804 => x"32700981",
   805 => x"05707207",
   806 => x"9f2a9171",
   807 => x"31515153",
   808 => x"53715183",
   809 => x"842d8114",
   810 => x"548e7425",
   811 => x"c23880c4",
   812 => x"f4085271",
   813 => x"80c6b40c",
   814 => x"0298050d",
   815 => x"0402f405",
   816 => x"0dd45281",
   817 => x"ff720c71",
   818 => x"085381ff",
   819 => x"720c7288",
   820 => x"2b83fe80",
   821 => x"06720870",
   822 => x"81ff0651",
   823 => x"525381ff",
   824 => x"720c7271",
   825 => x"07882b72",
   826 => x"087081ff",
   827 => x"06515253",
   828 => x"81ff720c",
   829 => x"72710788",
   830 => x"2b720870",
   831 => x"81ff0672",
   832 => x"0780c6b4",
   833 => x"0c525302",
   834 => x"8c050d04",
   835 => x"02f4050d",
   836 => x"74767181",
   837 => x"ff06d40c",
   838 => x"535380c7",
   839 => x"98088538",
   840 => x"71892b52",
   841 => x"71982ad4",
   842 => x"0c71902a",
   843 => x"7081ff06",
   844 => x"d40c5171",
   845 => x"882a7081",
   846 => x"ff06d40c",
   847 => x"517181ff",
   848 => x"06d40c72",
   849 => x"902a7081",
   850 => x"ff06d40c",
   851 => x"51d40870",
   852 => x"81ff0651",
   853 => x"5182b8bf",
   854 => x"527081ff",
   855 => x"2e098106",
   856 => x"943881ff",
   857 => x"0bd40cd4",
   858 => x"087081ff",
   859 => x"06ff1454",
   860 => x"515171e5",
   861 => x"387080c6",
   862 => x"b40c028c",
   863 => x"050d0402",
   864 => x"fc050d81",
   865 => x"c75181ff",
   866 => x"0bd40cff",
   867 => x"11517080",
   868 => x"25f43802",
   869 => x"84050d04",
   870 => x"02f4050d",
   871 => x"81ff0bd4",
   872 => x"0c935380",
   873 => x"5287fc80",
   874 => x"c1519a8c",
   875 => x"2d80c6b4",
   876 => x"088b3881",
   877 => x"ff0bd40c",
   878 => x"81539bc6",
   879 => x"049aff2d",
   880 => x"ff135372",
   881 => x"de387280",
   882 => x"c6b40c02",
   883 => x"8c050d04",
   884 => x"02ec050d",
   885 => x"810b80c7",
   886 => x"980c8454",
   887 => x"d008708f",
   888 => x"2a708106",
   889 => x"51515372",
   890 => x"f33872d0",
   891 => x"0c9aff2d",
   892 => x"bdd45186",
   893 => x"a02dd008",
   894 => x"708f2a70",
   895 => x"81065151",
   896 => x"5372f338",
   897 => x"810bd00c",
   898 => x"b1538052",
   899 => x"84d480c0",
   900 => x"519a8c2d",
   901 => x"80c6b408",
   902 => x"812e9338",
   903 => x"72822ebf",
   904 => x"38ff1353",
   905 => x"72e438ff",
   906 => x"145473ff",
   907 => x"af389aff",
   908 => x"2d83aa52",
   909 => x"849c80c8",
   910 => x"519a8c2d",
   911 => x"80c6b408",
   912 => x"812e0981",
   913 => x"06933899",
   914 => x"bd2d80c6",
   915 => x"b40883ff",
   916 => x"ff065372",
   917 => x"83aa2e9d",
   918 => x"389b982d",
   919 => x"9cf004bd",
   920 => x"e05186a0",
   921 => x"2d80539e",
   922 => x"c504bdf8",
   923 => x"5186a02d",
   924 => x"80549e96",
   925 => x"0481ff0b",
   926 => x"d40cb154",
   927 => x"9aff2d8f",
   928 => x"cf538052",
   929 => x"87fc80f7",
   930 => x"519a8c2d",
   931 => x"80c6b408",
   932 => x"5580c6b4",
   933 => x"08812e09",
   934 => x"81069c38",
   935 => x"81ff0bd4",
   936 => x"0c820a52",
   937 => x"849c80e9",
   938 => x"519a8c2d",
   939 => x"80c6b408",
   940 => x"802e8d38",
   941 => x"9aff2dff",
   942 => x"135372c6",
   943 => x"389e8904",
   944 => x"81ff0bd4",
   945 => x"0c80c6b4",
   946 => x"085287fc",
   947 => x"80fa519a",
   948 => x"8c2d80c6",
   949 => x"b408b238",
   950 => x"81ff0bd4",
   951 => x"0cd40853",
   952 => x"81ff0bd4",
   953 => x"0c81ff0b",
   954 => x"d40c81ff",
   955 => x"0bd40c81",
   956 => x"ff0bd40c",
   957 => x"72862a70",
   958 => x"81067656",
   959 => x"51537296",
   960 => x"3880c6b4",
   961 => x"08549e96",
   962 => x"0473822e",
   963 => x"fedc38ff",
   964 => x"145473fe",
   965 => x"e7387380",
   966 => x"c7980c73",
   967 => x"8b388152",
   968 => x"87fc80d0",
   969 => x"519a8c2d",
   970 => x"81ff0bd4",
   971 => x"0cd00870",
   972 => x"8f2a7081",
   973 => x"06515153",
   974 => x"72f33872",
   975 => x"d00c81ff",
   976 => x"0bd40c81",
   977 => x"537280c6",
   978 => x"b40c0294",
   979 => x"050d0402",
   980 => x"e8050d78",
   981 => x"55805681",
   982 => x"ff0bd40c",
   983 => x"d008708f",
   984 => x"2a708106",
   985 => x"51515372",
   986 => x"f3388281",
   987 => x"0bd00c81",
   988 => x"ff0bd40c",
   989 => x"775287fc",
   990 => x"80d1519a",
   991 => x"8c2d80db",
   992 => x"c6df5480",
   993 => x"c6b40880",
   994 => x"2e8a38be",
   995 => x"985186a0",
   996 => x"2d9fe804",
   997 => x"81ff0bd4",
   998 => x"0cd40870",
   999 => x"81ff0651",
  1000 => x"537281fe",
  1001 => x"2e098106",
  1002 => x"9e3880ff",
  1003 => x"5399bd2d",
  1004 => x"80c6b408",
  1005 => x"75708405",
  1006 => x"570cff13",
  1007 => x"53728025",
  1008 => x"ec388156",
  1009 => x"9fcd04ff",
  1010 => x"145473c8",
  1011 => x"3881ff0b",
  1012 => x"d40c81ff",
  1013 => x"0bd40cd0",
  1014 => x"08708f2a",
  1015 => x"70810651",
  1016 => x"515372f3",
  1017 => x"3872d00c",
  1018 => x"7580c6b4",
  1019 => x"0c029805",
  1020 => x"0d0402e8",
  1021 => x"050d7779",
  1022 => x"7b585555",
  1023 => x"80537276",
  1024 => x"25a33874",
  1025 => x"70810556",
  1026 => x"80f52d74",
  1027 => x"70810556",
  1028 => x"80f52d52",
  1029 => x"5271712e",
  1030 => x"86388151",
  1031 => x"a0a70481",
  1032 => x"13539ffe",
  1033 => x"04805170",
  1034 => x"80c6b40c",
  1035 => x"0298050d",
  1036 => x"0402ec05",
  1037 => x"0d765574",
  1038 => x"802e80c2",
  1039 => x"389a1580",
  1040 => x"e02d51ae",
  1041 => x"be2d80c6",
  1042 => x"b40880c6",
  1043 => x"b40880cd",
  1044 => x"cc0c80c6",
  1045 => x"b4085454",
  1046 => x"80cda808",
  1047 => x"802e9a38",
  1048 => x"941580e0",
  1049 => x"2d51aebe",
  1050 => x"2d80c6b4",
  1051 => x"08902b83",
  1052 => x"fff00a06",
  1053 => x"70750751",
  1054 => x"537280cd",
  1055 => x"cc0c80cd",
  1056 => x"cc085372",
  1057 => x"802e9d38",
  1058 => x"80cda008",
  1059 => x"fe147129",
  1060 => x"80cdb408",
  1061 => x"0580cdd0",
  1062 => x"0c70842b",
  1063 => x"80cdac0c",
  1064 => x"54a1d204",
  1065 => x"80cdb808",
  1066 => x"80cdcc0c",
  1067 => x"80cdbc08",
  1068 => x"80cdd00c",
  1069 => x"80cda808",
  1070 => x"802e8b38",
  1071 => x"80cda008",
  1072 => x"842b53a1",
  1073 => x"cd0480cd",
  1074 => x"c008842b",
  1075 => x"537280cd",
  1076 => x"ac0c0294",
  1077 => x"050d0402",
  1078 => x"d8050d80",
  1079 => x"0b80cda8",
  1080 => x"0c84549b",
  1081 => x"d02d80c6",
  1082 => x"b408802e",
  1083 => x"973880c7",
  1084 => x"9c528051",
  1085 => x"9ecf2d80",
  1086 => x"c6b40880",
  1087 => x"2e8638fe",
  1088 => x"54a28c04",
  1089 => x"ff145473",
  1090 => x"8024d838",
  1091 => x"738c38be",
  1092 => x"a85186a0",
  1093 => x"2d7355a7",
  1094 => x"d9048056",
  1095 => x"810b80cd",
  1096 => x"d40c8853",
  1097 => x"bebc5280",
  1098 => x"c7d2519f",
  1099 => x"f22d80c6",
  1100 => x"b408762e",
  1101 => x"09810689",
  1102 => x"3880c6b4",
  1103 => x"0880cdd4",
  1104 => x"0c8853be",
  1105 => x"c85280c7",
  1106 => x"ee519ff2",
  1107 => x"2d80c6b4",
  1108 => x"08893880",
  1109 => x"c6b40880",
  1110 => x"cdd40c80",
  1111 => x"cdd40880",
  1112 => x"2e818038",
  1113 => x"80cae20b",
  1114 => x"80f52d80",
  1115 => x"cae30b80",
  1116 => x"f52d7198",
  1117 => x"2b71902b",
  1118 => x"0780cae4",
  1119 => x"0b80f52d",
  1120 => x"70882b72",
  1121 => x"0780cae5",
  1122 => x"0b80f52d",
  1123 => x"710780cb",
  1124 => x"9a0b80f5",
  1125 => x"2d80cb9b",
  1126 => x"0b80f52d",
  1127 => x"71882b07",
  1128 => x"535f5452",
  1129 => x"5a565755",
  1130 => x"7381abaa",
  1131 => x"2e098106",
  1132 => x"8e387551",
  1133 => x"ae8d2d80",
  1134 => x"c6b40856",
  1135 => x"a3cc0473",
  1136 => x"82d4d52e",
  1137 => x"8738bed4",
  1138 => x"51a49504",
  1139 => x"80c79c52",
  1140 => x"75519ecf",
  1141 => x"2d80c6b4",
  1142 => x"085580c6",
  1143 => x"b408802e",
  1144 => x"83f73888",
  1145 => x"53bec852",
  1146 => x"80c7ee51",
  1147 => x"9ff22d80",
  1148 => x"c6b4088a",
  1149 => x"38810b80",
  1150 => x"cda80ca4",
  1151 => x"9b048853",
  1152 => x"bebc5280",
  1153 => x"c7d2519f",
  1154 => x"f22d80c6",
  1155 => x"b408802e",
  1156 => x"8a38bee8",
  1157 => x"5186a02d",
  1158 => x"a4fa0480",
  1159 => x"cb9a0b80",
  1160 => x"f52d5473",
  1161 => x"80d52e09",
  1162 => x"810680ce",
  1163 => x"3880cb9b",
  1164 => x"0b80f52d",
  1165 => x"547381aa",
  1166 => x"2e098106",
  1167 => x"bd38800b",
  1168 => x"80c79c0b",
  1169 => x"80f52d56",
  1170 => x"547481e9",
  1171 => x"2e833881",
  1172 => x"547481eb",
  1173 => x"2e8c3880",
  1174 => x"5573752e",
  1175 => x"09810682",
  1176 => x"f83880c7",
  1177 => x"a70b80f5",
  1178 => x"2d55748e",
  1179 => x"3880c7a8",
  1180 => x"0b80f52d",
  1181 => x"5473822e",
  1182 => x"86388055",
  1183 => x"a7d90480",
  1184 => x"c7a90b80",
  1185 => x"f52d7080",
  1186 => x"cda00cff",
  1187 => x"0580cda4",
  1188 => x"0c80c7aa",
  1189 => x"0b80f52d",
  1190 => x"80c7ab0b",
  1191 => x"80f52d58",
  1192 => x"76057782",
  1193 => x"80290570",
  1194 => x"80cdb00c",
  1195 => x"80c7ac0b",
  1196 => x"80f52d70",
  1197 => x"80cdc40c",
  1198 => x"80cda808",
  1199 => x"59575876",
  1200 => x"802e81b6",
  1201 => x"388853be",
  1202 => x"c85280c7",
  1203 => x"ee519ff2",
  1204 => x"2d80c6b4",
  1205 => x"08828238",
  1206 => x"80cda008",
  1207 => x"70842b80",
  1208 => x"cdac0c70",
  1209 => x"80cdc00c",
  1210 => x"80c7c10b",
  1211 => x"80f52d80",
  1212 => x"c7c00b80",
  1213 => x"f52d7182",
  1214 => x"80290580",
  1215 => x"c7c20b80",
  1216 => x"f52d7084",
  1217 => x"80802912",
  1218 => x"80c7c30b",
  1219 => x"80f52d70",
  1220 => x"81800a29",
  1221 => x"127080cd",
  1222 => x"c80c80cd",
  1223 => x"c4087129",
  1224 => x"80cdb008",
  1225 => x"057080cd",
  1226 => x"b40c80c7",
  1227 => x"c90b80f5",
  1228 => x"2d80c7c8",
  1229 => x"0b80f52d",
  1230 => x"71828029",
  1231 => x"0580c7ca",
  1232 => x"0b80f52d",
  1233 => x"70848080",
  1234 => x"291280c7",
  1235 => x"cb0b80f5",
  1236 => x"2d70982b",
  1237 => x"81f00a06",
  1238 => x"72057080",
  1239 => x"cdb80cfe",
  1240 => x"117e2977",
  1241 => x"0580cdbc",
  1242 => x"0c525952",
  1243 => x"43545e51",
  1244 => x"5259525d",
  1245 => x"575957a7",
  1246 => x"d20480c7",
  1247 => x"ae0b80f5",
  1248 => x"2d80c7ad",
  1249 => x"0b80f52d",
  1250 => x"71828029",
  1251 => x"057080cd",
  1252 => x"ac0c70a0",
  1253 => x"2983ff05",
  1254 => x"70892a70",
  1255 => x"80cdc00c",
  1256 => x"80c7b30b",
  1257 => x"80f52d80",
  1258 => x"c7b20b80",
  1259 => x"f52d7182",
  1260 => x"80290570",
  1261 => x"80cdc80c",
  1262 => x"7b71291e",
  1263 => x"7080cdbc",
  1264 => x"0c7d80cd",
  1265 => x"b80c7305",
  1266 => x"80cdb40c",
  1267 => x"555e5151",
  1268 => x"55558051",
  1269 => x"a0b12d81",
  1270 => x"557480c6",
  1271 => x"b40c02a8",
  1272 => x"050d0402",
  1273 => x"ec050d76",
  1274 => x"70872c71",
  1275 => x"80ff0655",
  1276 => x"565480cd",
  1277 => x"a8088a38",
  1278 => x"73882c74",
  1279 => x"81ff0654",
  1280 => x"5580c79c",
  1281 => x"5280cdb0",
  1282 => x"0815519e",
  1283 => x"cf2d80c6",
  1284 => x"b4085480",
  1285 => x"c6b40880",
  1286 => x"2eb83880",
  1287 => x"cda80880",
  1288 => x"2e9a3872",
  1289 => x"842980c7",
  1290 => x"9c057008",
  1291 => x"5253ae8d",
  1292 => x"2d80c6b4",
  1293 => x"08f00a06",
  1294 => x"53a8d004",
  1295 => x"721080c7",
  1296 => x"9c057080",
  1297 => x"e02d5253",
  1298 => x"aebe2d80",
  1299 => x"c6b40853",
  1300 => x"72547380",
  1301 => x"c6b40c02",
  1302 => x"94050d04",
  1303 => x"02e0050d",
  1304 => x"7970842c",
  1305 => x"80cdd008",
  1306 => x"05718f06",
  1307 => x"52555372",
  1308 => x"8a3880c7",
  1309 => x"9c527351",
  1310 => x"9ecf2d72",
  1311 => x"a02980c7",
  1312 => x"9c055480",
  1313 => x"7480f52d",
  1314 => x"56537473",
  1315 => x"2e833881",
  1316 => x"537481e5",
  1317 => x"2e81f438",
  1318 => x"81707406",
  1319 => x"54587280",
  1320 => x"2e81e838",
  1321 => x"8b1480f5",
  1322 => x"2d70832a",
  1323 => x"79065856",
  1324 => x"769b3880",
  1325 => x"c4f80853",
  1326 => x"72893872",
  1327 => x"80cb9c0b",
  1328 => x"81b72d76",
  1329 => x"80c4f80c",
  1330 => x"7353ab8d",
  1331 => x"04758f2e",
  1332 => x"09810681",
  1333 => x"b638749f",
  1334 => x"068d2980",
  1335 => x"cb8f1151",
  1336 => x"53811480",
  1337 => x"f52d7370",
  1338 => x"81055581",
  1339 => x"b72d8314",
  1340 => x"80f52d73",
  1341 => x"70810555",
  1342 => x"81b72d85",
  1343 => x"1480f52d",
  1344 => x"73708105",
  1345 => x"5581b72d",
  1346 => x"871480f5",
  1347 => x"2d737081",
  1348 => x"055581b7",
  1349 => x"2d891480",
  1350 => x"f52d7370",
  1351 => x"81055581",
  1352 => x"b72d8e14",
  1353 => x"80f52d73",
  1354 => x"70810555",
  1355 => x"81b72d90",
  1356 => x"1480f52d",
  1357 => x"73708105",
  1358 => x"5581b72d",
  1359 => x"921480f5",
  1360 => x"2d737081",
  1361 => x"055581b7",
  1362 => x"2d941480",
  1363 => x"f52d7370",
  1364 => x"81055581",
  1365 => x"b72d9614",
  1366 => x"80f52d73",
  1367 => x"70810555",
  1368 => x"81b72d98",
  1369 => x"1480f52d",
  1370 => x"73708105",
  1371 => x"5581b72d",
  1372 => x"9c1480f5",
  1373 => x"2d737081",
  1374 => x"055581b7",
  1375 => x"2d9e1480",
  1376 => x"f52d7381",
  1377 => x"b72d7780",
  1378 => x"c4f80c80",
  1379 => x"537280c6",
  1380 => x"b40c02a0",
  1381 => x"050d0402",
  1382 => x"cc050d7e",
  1383 => x"605e5a80",
  1384 => x"0b80cdcc",
  1385 => x"0880cdd0",
  1386 => x"08595c56",
  1387 => x"805880cd",
  1388 => x"ac08782e",
  1389 => x"81b83877",
  1390 => x"8f06a017",
  1391 => x"57547391",
  1392 => x"3880c79c",
  1393 => x"52765181",
  1394 => x"17579ecf",
  1395 => x"2d80c79c",
  1396 => x"56807680",
  1397 => x"f52d5654",
  1398 => x"74742e83",
  1399 => x"38815474",
  1400 => x"81e52e80",
  1401 => x"fd388170",
  1402 => x"7506555c",
  1403 => x"73802e80",
  1404 => x"f1388b16",
  1405 => x"80f52d98",
  1406 => x"06597880",
  1407 => x"e5388b53",
  1408 => x"7c527551",
  1409 => x"9ff22d80",
  1410 => x"c6b40880",
  1411 => x"d5389c16",
  1412 => x"0851ae8d",
  1413 => x"2d80c6b4",
  1414 => x"08841b0c",
  1415 => x"9a1680e0",
  1416 => x"2d51aebe",
  1417 => x"2d80c6b4",
  1418 => x"0880c6b4",
  1419 => x"08881c0c",
  1420 => x"80c6b408",
  1421 => x"555580cd",
  1422 => x"a808802e",
  1423 => x"99389416",
  1424 => x"80e02d51",
  1425 => x"aebe2d80",
  1426 => x"c6b40890",
  1427 => x"2b83fff0",
  1428 => x"0a067016",
  1429 => x"51547388",
  1430 => x"1b0c787a",
  1431 => x"0c7b54ad",
  1432 => x"aa048118",
  1433 => x"5880cdac",
  1434 => x"087826fe",
  1435 => x"ca3880cd",
  1436 => x"a808802e",
  1437 => x"b3387a51",
  1438 => x"a7e32d80",
  1439 => x"c6b40880",
  1440 => x"c6b40880",
  1441 => x"fffffff8",
  1442 => x"06555b73",
  1443 => x"80ffffff",
  1444 => x"f82e9538",
  1445 => x"80c6b408",
  1446 => x"fe0580cd",
  1447 => x"a0082980",
  1448 => x"cdb40805",
  1449 => x"57abac04",
  1450 => x"80547380",
  1451 => x"c6b40c02",
  1452 => x"b4050d04",
  1453 => x"02f4050d",
  1454 => x"74700881",
  1455 => x"05710c70",
  1456 => x"0880cda4",
  1457 => x"08065353",
  1458 => x"718f3888",
  1459 => x"130851a7",
  1460 => x"e32d80c6",
  1461 => x"b4088814",
  1462 => x"0c810b80",
  1463 => x"c6b40c02",
  1464 => x"8c050d04",
  1465 => x"02f0050d",
  1466 => x"75881108",
  1467 => x"fe0580cd",
  1468 => x"a0082980",
  1469 => x"cdb40811",
  1470 => x"720880cd",
  1471 => x"a4080605",
  1472 => x"79555354",
  1473 => x"549ecf2d",
  1474 => x"0290050d",
  1475 => x"0402f405",
  1476 => x"0d747088",
  1477 => x"2a83fe80",
  1478 => x"06707298",
  1479 => x"2a077288",
  1480 => x"2b87fc80",
  1481 => x"80067398",
  1482 => x"2b81f00a",
  1483 => x"06717307",
  1484 => x"0780c6b4",
  1485 => x"0c565153",
  1486 => x"51028c05",
  1487 => x"0d0402f8",
  1488 => x"050d028e",
  1489 => x"0580f52d",
  1490 => x"74882b07",
  1491 => x"7083ffff",
  1492 => x"0680c6b4",
  1493 => x"0c510288",
  1494 => x"050d0402",
  1495 => x"f4050d74",
  1496 => x"76785354",
  1497 => x"52807125",
  1498 => x"97387270",
  1499 => x"81055480",
  1500 => x"f52d7270",
  1501 => x"81055481",
  1502 => x"b72dff11",
  1503 => x"5170eb38",
  1504 => x"807281b7",
  1505 => x"2d028c05",
  1506 => x"0d0402e8",
  1507 => x"050d7756",
  1508 => x"80705654",
  1509 => x"737624b6",
  1510 => x"3880cdac",
  1511 => x"08742eae",
  1512 => x"387351a8",
  1513 => x"dc2d80c6",
  1514 => x"b40880c6",
  1515 => x"b4080981",
  1516 => x"057080c6",
  1517 => x"b408079f",
  1518 => x"2a770581",
  1519 => x"17575753",
  1520 => x"53747624",
  1521 => x"893880cd",
  1522 => x"ac087426",
  1523 => x"d4387280",
  1524 => x"c6b40c02",
  1525 => x"98050d04",
  1526 => x"02f0050d",
  1527 => x"80c6b008",
  1528 => x"1651af8a",
  1529 => x"2d80c6b4",
  1530 => x"08802e9f",
  1531 => x"388b5380",
  1532 => x"c6b40852",
  1533 => x"80cb9c51",
  1534 => x"aedb2d80",
  1535 => x"cdd80854",
  1536 => x"73802e87",
  1537 => x"3880cb9c",
  1538 => x"51732d02",
  1539 => x"90050d04",
  1540 => x"02dc050d",
  1541 => x"80705a55",
  1542 => x"7480c6b0",
  1543 => x"0825b438",
  1544 => x"80cdac08",
  1545 => x"752eac38",
  1546 => x"7851a8dc",
  1547 => x"2d80c6b4",
  1548 => x"08098105",
  1549 => x"7080c6b4",
  1550 => x"08079f2a",
  1551 => x"7605811b",
  1552 => x"5b565474",
  1553 => x"80c6b008",
  1554 => x"25893880",
  1555 => x"cdac0879",
  1556 => x"26d63880",
  1557 => x"557880cd",
  1558 => x"ac082781",
  1559 => x"db387851",
  1560 => x"a8dc2d80",
  1561 => x"c6b40880",
  1562 => x"2e81ad38",
  1563 => x"80c6b408",
  1564 => x"8b0580f5",
  1565 => x"2d70842a",
  1566 => x"70810677",
  1567 => x"1078842b",
  1568 => x"80cb9c0b",
  1569 => x"80f52d5c",
  1570 => x"5c535155",
  1571 => x"5673802e",
  1572 => x"80cb3874",
  1573 => x"16822bb2",
  1574 => x"dc0b80c5",
  1575 => x"84120c54",
  1576 => x"77753110",
  1577 => x"80cddc11",
  1578 => x"55569074",
  1579 => x"70810556",
  1580 => x"81b72da0",
  1581 => x"7481b72d",
  1582 => x"7681ff06",
  1583 => x"81165854",
  1584 => x"73802e8a",
  1585 => x"389c5380",
  1586 => x"cb9c52b1",
  1587 => x"d5048b53",
  1588 => x"80c6b408",
  1589 => x"5280cdde",
  1590 => x"1651b290",
  1591 => x"04741682",
  1592 => x"2bafd80b",
  1593 => x"80c58412",
  1594 => x"0c547681",
  1595 => x"ff068116",
  1596 => x"58547380",
  1597 => x"2e8a389c",
  1598 => x"5380cb9c",
  1599 => x"52b28704",
  1600 => x"8b5380c6",
  1601 => x"b4085277",
  1602 => x"75311080",
  1603 => x"cddc0551",
  1604 => x"7655aedb",
  1605 => x"2db2ad04",
  1606 => x"74902975",
  1607 => x"31701080",
  1608 => x"cddc0551",
  1609 => x"5480c6b4",
  1610 => x"087481b7",
  1611 => x"2d811959",
  1612 => x"748b24a3",
  1613 => x"38b0d504",
  1614 => x"74902975",
  1615 => x"31701080",
  1616 => x"cddc058c",
  1617 => x"77315751",
  1618 => x"54807481",
  1619 => x"b72d9e14",
  1620 => x"ff165654",
  1621 => x"74f33802",
  1622 => x"a4050d04",
  1623 => x"02fc050d",
  1624 => x"80c6b008",
  1625 => x"1351af8a",
  1626 => x"2d80c6b4",
  1627 => x"08802e89",
  1628 => x"3880c6b4",
  1629 => x"0851a0b1",
  1630 => x"2d800b80",
  1631 => x"c6b00cb0",
  1632 => x"902d9198",
  1633 => x"2d028405",
  1634 => x"0d0402fc",
  1635 => x"050d7251",
  1636 => x"70fd2eb0",
  1637 => x"3870fd24",
  1638 => x"8a3870fc",
  1639 => x"2e80cc38",
  1640 => x"b3f50470",
  1641 => x"fe2eb738",
  1642 => x"70ff2e09",
  1643 => x"810680c5",
  1644 => x"3880c6b0",
  1645 => x"08517080",
  1646 => x"2ebb38ff",
  1647 => x"1180c6b0",
  1648 => x"0cb3f504",
  1649 => x"80c6b008",
  1650 => x"f0057080",
  1651 => x"c6b00c51",
  1652 => x"708025a1",
  1653 => x"38800b80",
  1654 => x"c6b00cb3",
  1655 => x"f50480c6",
  1656 => x"b0088105",
  1657 => x"80c6b00c",
  1658 => x"b3f50480",
  1659 => x"c6b00890",
  1660 => x"0580c6b0",
  1661 => x"0cb0902d",
  1662 => x"91982d02",
  1663 => x"84050d04",
  1664 => x"02fc050d",
  1665 => x"800b80c6",
  1666 => x"b00cb090",
  1667 => x"2d90a82d",
  1668 => x"80c6b408",
  1669 => x"80c6a00c",
  1670 => x"80c4fc51",
  1671 => x"92bb2d02",
  1672 => x"84050d04",
  1673 => x"7180cdd8",
  1674 => x"0c040000",
  1675 => x"00ffffff",
  1676 => x"ff00ffff",
  1677 => x"ffff00ff",
  1678 => x"ffffff00",
  1679 => x"45786974",
  1680 => x"00000000",
  1681 => x"506f7420",
  1682 => x"33263420",
  1683 => x"4a6f7920",
  1684 => x"32204469",
  1685 => x"73706172",
  1686 => x"6f20322f",
  1687 => x"33000000",
  1688 => x"506f7420",
  1689 => x"33263420",
  1690 => x"5261746f",
  1691 => x"6e000000",
  1692 => x"506f7420",
  1693 => x"33263420",
  1694 => x"50616464",
  1695 => x"6c657320",
  1696 => x"33263400",
  1697 => x"506f7420",
  1698 => x"31263220",
  1699 => x"4a6f7920",
  1700 => x"31204469",
  1701 => x"73706172",
  1702 => x"6f20322f",
  1703 => x"33000000",
  1704 => x"506f7420",
  1705 => x"31263220",
  1706 => x"5261746f",
  1707 => x"6e000000",
  1708 => x"506f7420",
  1709 => x"31263220",
  1710 => x"50616464",
  1711 => x"6c657320",
  1712 => x"31263200",
  1713 => x"50756572",
  1714 => x"746f2055",
  1715 => x"41525400",
  1716 => x"50756572",
  1717 => x"746f204a",
  1718 => x"6f797374",
  1719 => x"69636b73",
  1720 => x"00000000",
  1721 => x"4a6f7973",
  1722 => x"7469636b",
  1723 => x"73204e6f",
  1724 => x"726d616c",
  1725 => x"00000000",
  1726 => x"4a6f7973",
  1727 => x"7469636b",
  1728 => x"7320496e",
  1729 => x"74657263",
  1730 => x"616d6269",
  1731 => x"61646f73",
  1732 => x"00000000",
  1733 => x"44696769",
  1734 => x"6d617820",
  1735 => x"4e6f0000",
  1736 => x"44696769",
  1737 => x"6d617820",
  1738 => x"24444530",
  1739 => x"30000000",
  1740 => x"44696769",
  1741 => x"6d617820",
  1742 => x"24444630",
  1743 => x"30000000",
  1744 => x"4d657a63",
  1745 => x"6c612053",
  1746 => x"74657265",
  1747 => x"6f204e6f",
  1748 => x"00000000",
  1749 => x"4d657a63",
  1750 => x"6c612053",
  1751 => x"74657265",
  1752 => x"6f203235",
  1753 => x"25000000",
  1754 => x"4d657a63",
  1755 => x"6c612053",
  1756 => x"74657265",
  1757 => x"6f203530",
  1758 => x"25000000",
  1759 => x"4d657a63",
  1760 => x"6c612053",
  1761 => x"74657265",
  1762 => x"6f203130",
  1763 => x"30250000",
  1764 => x"45787061",
  1765 => x"6e73696f",
  1766 => x"6e206465",
  1767 => x"20536f6e",
  1768 => x"69646f20",
  1769 => x"4e6f0000",
  1770 => x"45787061",
  1771 => x"6e73696f",
  1772 => x"6e206465",
  1773 => x"20536f6e",
  1774 => x"69646f20",
  1775 => x"4f504c32",
  1776 => x"00000000",
  1777 => x"53494420",
  1778 => x"44657265",
  1779 => x"63686f20",
  1780 => x"41646472",
  1781 => x"20496775",
  1782 => x"616c0000",
  1783 => x"53494420",
  1784 => x"44657265",
  1785 => x"63686f20",
  1786 => x"41646472",
  1787 => x"20244434",
  1788 => x"32300000",
  1789 => x"53494420",
  1790 => x"44657265",
  1791 => x"63686f20",
  1792 => x"41646472",
  1793 => x"20244435",
  1794 => x"30300000",
  1795 => x"53494420",
  1796 => x"44657265",
  1797 => x"63686f20",
  1798 => x"36353831",
  1799 => x"00000000",
  1800 => x"53494420",
  1801 => x"44657265",
  1802 => x"63686f20",
  1803 => x"38353830",
  1804 => x"00000000",
  1805 => x"53494420",
  1806 => x"497a7175",
  1807 => x"69657264",
  1808 => x"6f203635",
  1809 => x"38310000",
  1810 => x"53494420",
  1811 => x"497a7175",
  1812 => x"69657264",
  1813 => x"6f203835",
  1814 => x"38300000",
  1815 => x"50616c65",
  1816 => x"74612043",
  1817 => x"36340000",
  1818 => x"50616c65",
  1819 => x"74612043",
  1820 => x"65506543",
  1821 => x"65526100",
  1822 => x"50616c65",
  1823 => x"74612050",
  1824 => x"6570746f",
  1825 => x"00000000",
  1826 => x"50616c65",
  1827 => x"74612043",
  1828 => x"6f6d756e",
  1829 => x"69747900",
  1830 => x"5363616e",
  1831 => x"646f7562",
  1832 => x"6c657220",
  1833 => x"4e696e67",
  1834 => x"756e6f00",
  1835 => x"5363616e",
  1836 => x"646f7562",
  1837 => x"6c657220",
  1838 => x"43525420",
  1839 => x"32352500",
  1840 => x"5363616e",
  1841 => x"646f7562",
  1842 => x"6c657220",
  1843 => x"43525420",
  1844 => x"35302500",
  1845 => x"5363616e",
  1846 => x"646f7562",
  1847 => x"6c657220",
  1848 => x"43525420",
  1849 => x"37352500",
  1850 => x"466f726d",
  1851 => x"61746f20",
  1852 => x"4f726967",
  1853 => x"696e616c",
  1854 => x"00000000",
  1855 => x"466f726d",
  1856 => x"61746f20",
  1857 => x"50616e74",
  1858 => x"616c6c61",
  1859 => x"20436f6d",
  1860 => x"706c6574",
  1861 => x"61000000",
  1862 => x"466f726d",
  1863 => x"61746f20",
  1864 => x"5b415243",
  1865 => x"315d0000",
  1866 => x"466f726d",
  1867 => x"61746f20",
  1868 => x"5b415243",
  1869 => x"325d0000",
  1870 => x"41737065",
  1871 => x"63746f20",
  1872 => x"4f726967",
  1873 => x"696e616c",
  1874 => x"00000000",
  1875 => x"41737065",
  1876 => x"63746f20",
  1877 => x"416e6368",
  1878 => x"6f000000",
  1879 => x"56696465",
  1880 => x"6f205041",
  1881 => x"4c000000",
  1882 => x"56696465",
  1883 => x"6f204e54",
  1884 => x"53430000",
  1885 => x"2020203d",
  1886 => x"20434f4d",
  1887 => x"4f444f52",
  1888 => x"45202036",
  1889 => x"34203d20",
  1890 => x"20200000",
  1891 => x"20202020",
  1892 => x"20204e65",
  1893 => x"75726f52",
  1894 => x"756c657a",
  1895 => x"20202020",
  1896 => x"20200000",
  1897 => x"20202020",
  1898 => x"20202020",
  1899 => x"20202020",
  1900 => x"20202020",
  1901 => x"20202020",
  1902 => x"20200000",
  1903 => x"52657365",
  1904 => x"74000000",
  1905 => x"52657365",
  1906 => x"74202620",
  1907 => x"536f6c74",
  1908 => x"61722043",
  1909 => x"61727475",
  1910 => x"63686f00",
  1911 => x"56696465",
  1912 => x"6f201000",
  1913 => x"41756469",
  1914 => x"6f201000",
  1915 => x"50756572",
  1916 => x"746f7320",
  1917 => x"10000000",
  1918 => x"53616361",
  1919 => x"72204369",
  1920 => x"6e746100",
  1921 => x"506c6179",
  1922 => x"2f53746f",
  1923 => x"70204369",
  1924 => x"6e746100",
  1925 => x"43617267",
  1926 => x"61722044",
  1927 => x"6973636f",
  1928 => x"2f43696e",
  1929 => x"74612f43",
  1930 => x"61727420",
  1931 => x"10000000",
  1932 => x"44697363",
  1933 => x"6f204772",
  1934 => x"61626162",
  1935 => x"6c650000",
  1936 => x"44697363",
  1937 => x"6f20536f",
  1938 => x"6c6f204c",
  1939 => x"65637475",
  1940 => x"72610000",
  1941 => x"536f6e69",
  1942 => x"646f2043",
  1943 => x"696e7461",
  1944 => x"204f6666",
  1945 => x"00000000",
  1946 => x"536f6e69",
  1947 => x"646f2043",
  1948 => x"696e7461",
  1949 => x"204f6e00",
  1950 => x"4b65726e",
  1951 => x"656c2043",
  1952 => x"61726761",
  1953 => x"626c6500",
  1954 => x"4b65726e",
  1955 => x"656c2043",
  1956 => x"36340000",
  1957 => x"4b65726e",
  1958 => x"656c2043",
  1959 => x"36344753",
  1960 => x"00000000",
  1961 => x"4b65726e",
  1962 => x"656c204a",
  1963 => x"61706f6e",
  1964 => x"65730000",
  1965 => x"43617267",
  1966 => x"61204661",
  1967 => x"6c6c6964",
  1968 => x"61000000",
  1969 => x"4f4b0000",
  1970 => x"16200000",
  1971 => x"14200000",
  1972 => x"15200000",
  1973 => x"53442069",
  1974 => x"6e69742e",
  1975 => x"2e2e0a00",
  1976 => x"53442063",
  1977 => x"61726420",
  1978 => x"72657365",
  1979 => x"74206661",
  1980 => x"696c6564",
  1981 => x"210a0000",
  1982 => x"53444843",
  1983 => x"20657272",
  1984 => x"6f72210a",
  1985 => x"00000000",
  1986 => x"57726974",
  1987 => x"65206661",
  1988 => x"696c6564",
  1989 => x"0a000000",
  1990 => x"52656164",
  1991 => x"20666169",
  1992 => x"6c65640a",
  1993 => x"00000000",
  1994 => x"43617264",
  1995 => x"20696e69",
  1996 => x"74206661",
  1997 => x"696c6564",
  1998 => x"0a000000",
  1999 => x"46415431",
  2000 => x"36202020",
  2001 => x"00000000",
  2002 => x"46415433",
  2003 => x"32202020",
  2004 => x"00000000",
  2005 => x"4e6f2070",
  2006 => x"61727469",
  2007 => x"74696f6e",
  2008 => x"20736967",
  2009 => x"0a000000",
  2010 => x"42616420",
  2011 => x"70617274",
  2012 => x"0a000000",
  2013 => x"4261636b",
  2014 => x"00000000",
  2015 => x"00000002",
  2016 => x"00000003",
  2017 => x"00001fe8",
  2018 => x"00000002",
  2019 => x"00000003",
  2020 => x"00001fe0",
  2021 => x"00000002",
  2022 => x"00000003",
  2023 => x"00001fd4",
  2024 => x"00000003",
  2025 => x"00000003",
  2026 => x"00001fc8",
  2027 => x"00000003",
  2028 => x"00000004",
  2029 => x"00001a3c",
  2030 => x"00002124",
  2031 => x"00000000",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00001a44",
  2035 => x"00001a60",
  2036 => x"00001a70",
  2037 => x"00001a84",
  2038 => x"00001aa0",
  2039 => x"00001ab0",
  2040 => x"00001ac4",
  2041 => x"00001ad0",
  2042 => x"00001ae4",
  2043 => x"00001af8",
  2044 => x"00000003",
  2045 => x"00002088",
  2046 => x"00000002",
  2047 => x"00000003",
  2048 => x"00002080",
  2049 => x"00000002",
  2050 => x"00000003",
  2051 => x"00002074",
  2052 => x"00000003",
  2053 => x"00000003",
  2054 => x"0000206c",
  2055 => x"00000002",
  2056 => x"00000003",
  2057 => x"0000205c",
  2058 => x"00000004",
  2059 => x"00000003",
  2060 => x"00002050",
  2061 => x"00000003",
  2062 => x"00000004",
  2063 => x"00001a3c",
  2064 => x"00002124",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00001b14",
  2069 => x"00001b20",
  2070 => x"00001b30",
  2071 => x"00001b40",
  2072 => x"00001b54",
  2073 => x"00001b68",
  2074 => x"00001b7c",
  2075 => x"00001b90",
  2076 => x"00001ba8",
  2077 => x"00001bc4",
  2078 => x"00001bdc",
  2079 => x"00001bf4",
  2080 => x"00001c0c",
  2081 => x"00001c20",
  2082 => x"00001c34",
  2083 => x"00001c48",
  2084 => x"00000003",
  2085 => x"0000211c",
  2086 => x"00000002",
  2087 => x"00000003",
  2088 => x"00002114",
  2089 => x"00000002",
  2090 => x"00000003",
  2091 => x"00002104",
  2092 => x"00000004",
  2093 => x"00000003",
  2094 => x"000020f4",
  2095 => x"00000004",
  2096 => x"00000003",
  2097 => x"000020e4",
  2098 => x"00000004",
  2099 => x"00000004",
  2100 => x"00001a3c",
  2101 => x"00002124",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00001c5c",
  2106 => x"00001c68",
  2107 => x"00001c78",
  2108 => x"00001c88",
  2109 => x"00001c98",
  2110 => x"00001cac",
  2111 => x"00001cc0",
  2112 => x"00001cd4",
  2113 => x"00001ce8",
  2114 => x"00001cfc",
  2115 => x"00001d18",
  2116 => x"00001d28",
  2117 => x"00001d38",
  2118 => x"00001d4c",
  2119 => x"00001d5c",
  2120 => x"00001d68",
  2121 => x"00000002",
  2122 => x"00001d74",
  2123 => x"00000000",
  2124 => x"00000002",
  2125 => x"00001d8c",
  2126 => x"00000000",
  2127 => x"00000002",
  2128 => x"00001da4",
  2129 => x"00000000",
  2130 => x"00000002",
  2131 => x"00001dbc",
  2132 => x"00000371",
  2133 => x"00000002",
  2134 => x"00001dc4",
  2135 => x"00000388",
  2136 => x"00000004",
  2137 => x"00001ddc",
  2138 => x"00002090",
  2139 => x"00000004",
  2140 => x"00001de4",
  2141 => x"00001ff0",
  2142 => x"00000004",
  2143 => x"00001dec",
  2144 => x"00001f80",
  2145 => x"00000003",
  2146 => x"000021f4",
  2147 => x"00000004",
  2148 => x"00000003",
  2149 => x"000021ec",
  2150 => x"00000002",
  2151 => x"00000003",
  2152 => x"000021e4",
  2153 => x"00000002",
  2154 => x"00000002",
  2155 => x"00001df8",
  2156 => x"000003b8",
  2157 => x"00000002",
  2158 => x"00001e04",
  2159 => x"000003a0",
  2160 => x"00000002",
  2161 => x"00001e14",
  2162 => x"00001a00",
  2163 => x"00000002",
  2164 => x"00001a3c",
  2165 => x"00000831",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00001e30",
  2170 => x"00001e40",
  2171 => x"00001e54",
  2172 => x"00001e68",
  2173 => x"00001e78",
  2174 => x"00001e88",
  2175 => x"00001e94",
  2176 => x"00001ea4",
  2177 => x"00000004",
  2178 => x"00001eb4",
  2179 => x"00002204",
  2180 => x"00000004",
  2181 => x"00001ec4",
  2182 => x"00002124",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000002",
  2208 => x"000026dc",
  2209 => x"000017d8",
  2210 => x"00000002",
  2211 => x"000026fa",
  2212 => x"000017d8",
  2213 => x"00000002",
  2214 => x"00002718",
  2215 => x"000017d8",
  2216 => x"00000002",
  2217 => x"00002736",
  2218 => x"000017d8",
  2219 => x"00000002",
  2220 => x"00002754",
  2221 => x"000017d8",
  2222 => x"00000002",
  2223 => x"00002772",
  2224 => x"000017d8",
  2225 => x"00000002",
  2226 => x"00002790",
  2227 => x"000017d8",
  2228 => x"00000002",
  2229 => x"000027ae",
  2230 => x"000017d8",
  2231 => x"00000002",
  2232 => x"000027cc",
  2233 => x"000017d8",
  2234 => x"00000002",
  2235 => x"000027ea",
  2236 => x"000017d8",
  2237 => x"00000002",
  2238 => x"00002808",
  2239 => x"000017d8",
  2240 => x"00000002",
  2241 => x"00002826",
  2242 => x"000017d8",
  2243 => x"00000002",
  2244 => x"00002844",
  2245 => x"000017d8",
  2246 => x"00000004",
  2247 => x"00001f74",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"0000198a",
  2252 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

