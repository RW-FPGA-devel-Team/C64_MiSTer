-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c6",
     9 => x"94080b0b",
    10 => x"80c69808",
    11 => x"0b0b80c6",
    12 => x"9c080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c69c0c0b",
    16 => x"0b80c698",
    17 => x"0c0b0b80",
    18 => x"c6940c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb49c",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c69470",
    57 => x"80d0c427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5189dd",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c6",
    65 => x"a40c9f0b",
    66 => x"80c6a80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c6a808ff",
    70 => x"0580c6a8",
    71 => x"0c80c6a8",
    72 => x"088025e8",
    73 => x"3880c6a4",
    74 => x"08ff0580",
    75 => x"c6a40c80",
    76 => x"c6a40880",
    77 => x"25d03880",
    78 => x"0b80c6a8",
    79 => x"0c800b80",
    80 => x"c6a40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c6a408",
   100 => x"25913882",
   101 => x"c82d80c6",
   102 => x"a408ff05",
   103 => x"80c6a40c",
   104 => x"838a0480",
   105 => x"c6a40880",
   106 => x"c6a80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c6a408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c6a80881",
   116 => x"0580c6a8",
   117 => x"0c80c6a8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c6a8",
   121 => x"0c80c6a4",
   122 => x"08810580",
   123 => x"c6a40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c6",
   128 => x"a8088105",
   129 => x"80c6a80c",
   130 => x"80c6a808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c6a8",
   134 => x"0c80c6a4",
   135 => x"08810580",
   136 => x"c6a40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"c6ac0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"c6ac0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280c6",
   177 => x"ac088407",
   178 => x"80c6ac0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b0bbe",
   183 => x"f00c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80c6ac",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80c6",
   208 => x"940c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050d84bf",
   216 => x"5186c72d",
   217 => x"ff115170",
   218 => x"8025f638",
   219 => x"0284050d",
   220 => x"0402fc05",
   221 => x"0dec5183",
   222 => x"710c86c7",
   223 => x"2d82710c",
   224 => x"90a22d02",
   225 => x"84050d04",
   226 => x"02fc050d",
   227 => x"ec518182",
   228 => x"710c86c7",
   229 => x"2d82710c",
   230 => x"90a22d02",
   231 => x"84050d04",
   232 => x"02fc050d",
   233 => x"ec5180c2",
   234 => x"710c86c7",
   235 => x"2d82710c",
   236 => x"90a22d02",
   237 => x"84050d04",
   238 => x"02fc050d",
   239 => x"ec518282",
   240 => x"710c86c7",
   241 => x"2d82710c",
   242 => x"90a22d02",
   243 => x"84050d04",
   244 => x"02fc050d",
   245 => x"ec519271",
   246 => x"0c86c72d",
   247 => x"82710c02",
   248 => x"84050d04",
   249 => x"02d0050d",
   250 => x"7d548074",
   251 => x"5380c6b0",
   252 => x"525bab88",
   253 => x"2d80c694",
   254 => x"087b2e81",
   255 => x"b63880c6",
   256 => x"b40870f8",
   257 => x"0c891580",
   258 => x"f52d8a16",
   259 => x"80f52d71",
   260 => x"82802905",
   261 => x"881780f5",
   262 => x"2d708480",
   263 => x"802912f4",
   264 => x"0c575556",
   265 => x"58a40bec",
   266 => x"0c7aff19",
   267 => x"585a767b",
   268 => x"2e8b3881",
   269 => x"1a77812a",
   270 => x"585a76f7",
   271 => x"38f71a5a",
   272 => x"815b8078",
   273 => x"2580ec38",
   274 => x"79527651",
   275 => x"84a82d80",
   276 => x"c6fc5280",
   277 => x"c6b051ad",
   278 => x"d52d80c6",
   279 => x"9408802e",
   280 => x"b93880c6",
   281 => x"fc5c83fc",
   282 => x"597b7084",
   283 => x"055d0870",
   284 => x"81ff0671",
   285 => x"882a7081",
   286 => x"ff067390",
   287 => x"2a7081ff",
   288 => x"0675982a",
   289 => x"e80ce80c",
   290 => x"58e80c57",
   291 => x"e80cfc1a",
   292 => x"5a537880",
   293 => x"25d33889",
   294 => x"a20480c6",
   295 => x"94085b84",
   296 => x"805880c6",
   297 => x"b051ada5",
   298 => x"2dfc8018",
   299 => x"81185858",
   300 => x"88c20486",
   301 => x"da2d840b",
   302 => x"ec0c7a80",
   303 => x"2e8e3880",
   304 => x"c2885192",
   305 => x"ac2d90a2",
   306 => x"2d89d304",
   307 => x"80c3e451",
   308 => x"92ac2d7a",
   309 => x"80c6940c",
   310 => x"02b0050d",
   311 => x"0402ec05",
   312 => x"0d840bec",
   313 => x"0c90802d",
   314 => x"8cd22d81",
   315 => x"f92da1c8",
   316 => x"2d80c694",
   317 => x"08802e82",
   318 => x"c23887e4",
   319 => x"51b4952d",
   320 => x"80c28851",
   321 => x"92ac2d90",
   322 => x"a22d8cde",
   323 => x"2d92bf2d",
   324 => x"80c1900b",
   325 => x"80f52d70",
   326 => x"822b8406",
   327 => x"80c19c0b",
   328 => x"80f52d70",
   329 => x"982b8180",
   330 => x"0a0680c1",
   331 => x"a80b80f5",
   332 => x"2d70842b",
   333 => x"b0067473",
   334 => x"070780c1",
   335 => x"b40b80f5",
   336 => x"2d70882b",
   337 => x"8e8006bf",
   338 => x"ec0b80f5",
   339 => x"2d708d2b",
   340 => x"80c08006",
   341 => x"74730707",
   342 => x"bff80b80",
   343 => x"f52d7090",
   344 => x"2b848080",
   345 => x"0680c084",
   346 => x"0b80f52d",
   347 => x"70942b9c",
   348 => x"800a0674",
   349 => x"73070780",
   350 => x"c0900b80",
   351 => x"f52d7086",
   352 => x"2b80c006",
   353 => x"80c09c0b",
   354 => x"80f52d70",
   355 => x"8c2ba080",
   356 => x"06747307",
   357 => x"0780c0a8",
   358 => x"0b80f52d",
   359 => x"70922bb0",
   360 => x"808006be",
   361 => x"fc0b80f5",
   362 => x"2d70832b",
   363 => x"88067473",
   364 => x"0707bf88",
   365 => x"0b80f52d",
   366 => x"70108206",
   367 => x"bf940b80",
   368 => x"f52d709a",
   369 => x"2bb00a06",
   370 => x"74730707",
   371 => x"bfa00b80",
   372 => x"f52d709c",
   373 => x"2b8c0a06",
   374 => x"80c2f00b",
   375 => x"80f52d70",
   376 => x"8e2b8380",
   377 => x"80067473",
   378 => x"070780c2",
   379 => x"fc0b80f5",
   380 => x"2d708b2b",
   381 => x"90800680",
   382 => x"c3880b80",
   383 => x"f52d709e",
   384 => x"2b820a06",
   385 => x"74730707",
   386 => x"fc0c5454",
   387 => x"54545454",
   388 => x"54545454",
   389 => x"54545454",
   390 => x"54545454",
   391 => x"54545454",
   392 => x"54545454",
   393 => x"56545257",
   394 => x"57535386",
   395 => x"5280c694",
   396 => x"08833884",
   397 => x"5271ec0c",
   398 => x"8a8a0480",
   399 => x"0b80c694",
   400 => x"0c029405",
   401 => x"0d047198",
   402 => x"0c04ffb0",
   403 => x"0880c694",
   404 => x"0c04810b",
   405 => x"ffb00c04",
   406 => x"800bffb0",
   407 => x"0c0402f4",
   408 => x"050d8dec",
   409 => x"0480c694",
   410 => x"0881f02e",
   411 => x"0981068a",
   412 => x"38810b80",
   413 => x"c4c80c8d",
   414 => x"ec0480c6",
   415 => x"940881e0",
   416 => x"2e098106",
   417 => x"8a38810b",
   418 => x"80c4cc0c",
   419 => x"8dec0480",
   420 => x"c6940852",
   421 => x"80c4cc08",
   422 => x"802e8938",
   423 => x"80c69408",
   424 => x"81800552",
   425 => x"71842c72",
   426 => x"8f065353",
   427 => x"80c4c808",
   428 => x"802e9a38",
   429 => x"72842980",
   430 => x"c4880572",
   431 => x"1381712b",
   432 => x"70097308",
   433 => x"06730c51",
   434 => x"53538de0",
   435 => x"04728429",
   436 => x"80c48805",
   437 => x"72138371",
   438 => x"2b720807",
   439 => x"720c5353",
   440 => x"800b80c4",
   441 => x"cc0c800b",
   442 => x"80c4c80c",
   443 => x"80c6bc51",
   444 => x"8ef32d80",
   445 => x"c69408ff",
   446 => x"24feea38",
   447 => x"800b80c6",
   448 => x"940c028c",
   449 => x"050d0402",
   450 => x"f8050d80",
   451 => x"c488528f",
   452 => x"51807270",
   453 => x"8405540c",
   454 => x"ff115170",
   455 => x"8025f238",
   456 => x"0288050d",
   457 => x"0402f005",
   458 => x"0d75518c",
   459 => x"d82d7082",
   460 => x"2cfc0680",
   461 => x"c4881172",
   462 => x"109e0671",
   463 => x"0870722a",
   464 => x"70830682",
   465 => x"742b7009",
   466 => x"7406760c",
   467 => x"54515657",
   468 => x"5351538c",
   469 => x"d22d7180",
   470 => x"c6940c02",
   471 => x"90050d04",
   472 => x"02fc050d",
   473 => x"72518071",
   474 => x"0c800b84",
   475 => x"120c0284",
   476 => x"050d0402",
   477 => x"f0050d75",
   478 => x"70088412",
   479 => x"08535353",
   480 => x"ff547171",
   481 => x"2ea8388c",
   482 => x"d82d8413",
   483 => x"08708429",
   484 => x"14881170",
   485 => x"087081ff",
   486 => x"06841808",
   487 => x"81118706",
   488 => x"841a0c53",
   489 => x"51555151",
   490 => x"518cd22d",
   491 => x"71547380",
   492 => x"c6940c02",
   493 => x"90050d04",
   494 => x"02f8050d",
   495 => x"8cd82de0",
   496 => x"08708b2a",
   497 => x"70810651",
   498 => x"52527080",
   499 => x"2ea13880",
   500 => x"c6bc0870",
   501 => x"842980c6",
   502 => x"c4057381",
   503 => x"ff06710c",
   504 => x"515180c6",
   505 => x"bc088111",
   506 => x"870680c6",
   507 => x"bc0c5180",
   508 => x"0b80c6e4",
   509 => x"0c8cca2d",
   510 => x"8cd22d02",
   511 => x"88050d04",
   512 => x"02fc050d",
   513 => x"80c6bc51",
   514 => x"8ee02d8e",
   515 => x"872d8fb8",
   516 => x"518cc62d",
   517 => x"0284050d",
   518 => x"0480c6e8",
   519 => x"0880c694",
   520 => x"0c0402fc",
   521 => x"050d90ac",
   522 => x"048cde2d",
   523 => x"80f6518e",
   524 => x"a52d80c6",
   525 => x"9408f238",
   526 => x"80da518e",
   527 => x"a52d80c6",
   528 => x"9408e638",
   529 => x"80c69408",
   530 => x"80c4d40c",
   531 => x"80c69408",
   532 => x"51858d2d",
   533 => x"0284050d",
   534 => x"0402ec05",
   535 => x"0d765480",
   536 => x"52870b88",
   537 => x"1580f52d",
   538 => x"56537472",
   539 => x"248338a0",
   540 => x"53725183",
   541 => x"842d8112",
   542 => x"8b1580f5",
   543 => x"2d545272",
   544 => x"7225de38",
   545 => x"0294050d",
   546 => x"0402f005",
   547 => x"0d80c6e8",
   548 => x"085481f9",
   549 => x"2d800b80",
   550 => x"c6ec0c73",
   551 => x"08802e81",
   552 => x"8638820b",
   553 => x"80c6a80c",
   554 => x"80c6ec08",
   555 => x"8f0680c6",
   556 => x"a40c7308",
   557 => x"5271832e",
   558 => x"96387183",
   559 => x"26893871",
   560 => x"812eaf38",
   561 => x"92900471",
   562 => x"852e9f38",
   563 => x"92900488",
   564 => x"1480f52d",
   565 => x"841508bd",
   566 => x"bc535452",
   567 => x"86a02d71",
   568 => x"84291370",
   569 => x"08525292",
   570 => x"94047351",
   571 => x"90d92d92",
   572 => x"900480c4",
   573 => x"d0088815",
   574 => x"082c7081",
   575 => x"06515271",
   576 => x"802e8738",
   577 => x"bdc05192",
   578 => x"8d04bdc4",
   579 => x"5186a02d",
   580 => x"84140851",
   581 => x"86a02d80",
   582 => x"c6ec0881",
   583 => x"0580c6ec",
   584 => x"0c8c1454",
   585 => x"919b0402",
   586 => x"90050d04",
   587 => x"7180c6e8",
   588 => x"0c91892d",
   589 => x"80c6ec08",
   590 => x"ff0580c6",
   591 => x"f00c0402",
   592 => x"e8050d80",
   593 => x"c6e80880",
   594 => x"c6f40857",
   595 => x"5587518e",
   596 => x"a52d80c6",
   597 => x"9408812a",
   598 => x"70810651",
   599 => x"5271802e",
   600 => x"a33892e8",
   601 => x"048cde2d",
   602 => x"87518ea5",
   603 => x"2d80c694",
   604 => x"08f33880",
   605 => x"c4d40881",
   606 => x"327080c4",
   607 => x"d40c7052",
   608 => x"52858d2d",
   609 => x"80fe518e",
   610 => x"a52d80c6",
   611 => x"9408802e",
   612 => x"a93880c4",
   613 => x"d408802e",
   614 => x"9238800b",
   615 => x"80c4d40c",
   616 => x"8051858d",
   617 => x"2d93ab04",
   618 => x"8cde2d80",
   619 => x"fe518ea5",
   620 => x"2d80c694",
   621 => x"08f23887",
   622 => x"d02d80c4",
   623 => x"d4089038",
   624 => x"81fd518e",
   625 => x"a52d81fa",
   626 => x"518ea52d",
   627 => x"99a40481",
   628 => x"f5518ea5",
   629 => x"2d80c694",
   630 => x"08812a70",
   631 => x"81065152",
   632 => x"71802eb3",
   633 => x"3880c6f0",
   634 => x"08527180",
   635 => x"2e8a38ff",
   636 => x"1280c6f0",
   637 => x"0c949704",
   638 => x"80c6ec08",
   639 => x"1080c6ec",
   640 => x"08057084",
   641 => x"29165152",
   642 => x"88120880",
   643 => x"2e8938ff",
   644 => x"51881208",
   645 => x"52712d81",
   646 => x"f2518ea5",
   647 => x"2d80c694",
   648 => x"08812a70",
   649 => x"81065152",
   650 => x"71802eb4",
   651 => x"3880c6ec",
   652 => x"08ff1180",
   653 => x"c6f00856",
   654 => x"53537372",
   655 => x"258a3881",
   656 => x"1480c6f0",
   657 => x"0c94e004",
   658 => x"72101370",
   659 => x"84291651",
   660 => x"52881208",
   661 => x"802e8938",
   662 => x"fe518812",
   663 => x"0852712d",
   664 => x"81fd518e",
   665 => x"a52d80c6",
   666 => x"9408812a",
   667 => x"70810651",
   668 => x"5271802e",
   669 => x"b13880c6",
   670 => x"f008802e",
   671 => x"8a38800b",
   672 => x"80c6f00c",
   673 => x"95a60480",
   674 => x"c6ec0810",
   675 => x"80c6ec08",
   676 => x"05708429",
   677 => x"16515288",
   678 => x"1208802e",
   679 => x"8938fd51",
   680 => x"88120852",
   681 => x"712d81fa",
   682 => x"518ea52d",
   683 => x"80c69408",
   684 => x"812a7081",
   685 => x"06515271",
   686 => x"802eb138",
   687 => x"80c6ec08",
   688 => x"ff115452",
   689 => x"80c6f008",
   690 => x"73258938",
   691 => x"7280c6f0",
   692 => x"0c95ec04",
   693 => x"71101270",
   694 => x"84291651",
   695 => x"52881208",
   696 => x"802e8938",
   697 => x"fc518812",
   698 => x"0852712d",
   699 => x"80c6f008",
   700 => x"70535473",
   701 => x"802e8a38",
   702 => x"8c15ff15",
   703 => x"555595f3",
   704 => x"04820b80",
   705 => x"c6a80c71",
   706 => x"8f0680c6",
   707 => x"a40c81eb",
   708 => x"518ea52d",
   709 => x"80c69408",
   710 => x"812a7081",
   711 => x"06515271",
   712 => x"802ead38",
   713 => x"7408852e",
   714 => x"098106a4",
   715 => x"38881580",
   716 => x"f52dff05",
   717 => x"52718816",
   718 => x"81b72d71",
   719 => x"982b5271",
   720 => x"80258838",
   721 => x"800b8816",
   722 => x"81b72d74",
   723 => x"5190d92d",
   724 => x"81f4518e",
   725 => x"a52d80c6",
   726 => x"9408812a",
   727 => x"70810651",
   728 => x"5271802e",
   729 => x"b3387408",
   730 => x"852e0981",
   731 => x"06aa3888",
   732 => x"1580f52d",
   733 => x"81055271",
   734 => x"881681b7",
   735 => x"2d7181ff",
   736 => x"068b1680",
   737 => x"f52d5452",
   738 => x"72722787",
   739 => x"38728816",
   740 => x"81b72d74",
   741 => x"5190d92d",
   742 => x"80da518e",
   743 => x"a52d80c6",
   744 => x"9408812a",
   745 => x"70810651",
   746 => x"5271802e",
   747 => x"81ad3880",
   748 => x"c6e80880",
   749 => x"c6f00855",
   750 => x"5373802e",
   751 => x"8a388c13",
   752 => x"ff155553",
   753 => x"97b90472",
   754 => x"08527182",
   755 => x"2ea63871",
   756 => x"82268938",
   757 => x"71812eaa",
   758 => x"3898db04",
   759 => x"71832eb4",
   760 => x"3871842e",
   761 => x"09810680",
   762 => x"f2388813",
   763 => x"085192ac",
   764 => x"2d98db04",
   765 => x"80c6f008",
   766 => x"51881308",
   767 => x"52712d98",
   768 => x"db04810b",
   769 => x"8814082b",
   770 => x"80c4d008",
   771 => x"3280c4d0",
   772 => x"0c98af04",
   773 => x"881380f5",
   774 => x"2d81058b",
   775 => x"1480f52d",
   776 => x"53547174",
   777 => x"24833880",
   778 => x"54738814",
   779 => x"81b72d91",
   780 => x"892d98db",
   781 => x"04750880",
   782 => x"2ea43875",
   783 => x"08518ea5",
   784 => x"2d80c694",
   785 => x"08810652",
   786 => x"71802e8c",
   787 => x"3880c6f0",
   788 => x"08518416",
   789 => x"0852712d",
   790 => x"88165675",
   791 => x"d8388054",
   792 => x"800b80c6",
   793 => x"a80c738f",
   794 => x"0680c6a4",
   795 => x"0ca05273",
   796 => x"80c6f008",
   797 => x"2e098106",
   798 => x"993880c6",
   799 => x"ec08ff05",
   800 => x"74327009",
   801 => x"81057072",
   802 => x"079f2a91",
   803 => x"71315151",
   804 => x"53537151",
   805 => x"83842d81",
   806 => x"14548e74",
   807 => x"25c23880",
   808 => x"c4d40852",
   809 => x"7180c694",
   810 => x"0c029805",
   811 => x"0d0402f4",
   812 => x"050dd452",
   813 => x"81ff720c",
   814 => x"71085381",
   815 => x"ff720c72",
   816 => x"882b83fe",
   817 => x"80067208",
   818 => x"7081ff06",
   819 => x"51525381",
   820 => x"ff720c72",
   821 => x"7107882b",
   822 => x"72087081",
   823 => x"ff065152",
   824 => x"5381ff72",
   825 => x"0c727107",
   826 => x"882b7208",
   827 => x"7081ff06",
   828 => x"720780c6",
   829 => x"940c5253",
   830 => x"028c050d",
   831 => x"0402f405",
   832 => x"0d747671",
   833 => x"81ff06d4",
   834 => x"0c535380",
   835 => x"c6f80885",
   836 => x"3871892b",
   837 => x"5271982a",
   838 => x"d40c7190",
   839 => x"2a7081ff",
   840 => x"06d40c51",
   841 => x"71882a70",
   842 => x"81ff06d4",
   843 => x"0c517181",
   844 => x"ff06d40c",
   845 => x"72902a70",
   846 => x"81ff06d4",
   847 => x"0c51d408",
   848 => x"7081ff06",
   849 => x"515182b8",
   850 => x"bf527081",
   851 => x"ff2e0981",
   852 => x"06943881",
   853 => x"ff0bd40c",
   854 => x"d4087081",
   855 => x"ff06ff14",
   856 => x"54515171",
   857 => x"e5387080",
   858 => x"c6940c02",
   859 => x"8c050d04",
   860 => x"02fc050d",
   861 => x"81c75181",
   862 => x"ff0bd40c",
   863 => x"ff115170",
   864 => x"8025f438",
   865 => x"0284050d",
   866 => x"0402f405",
   867 => x"0d81ff0b",
   868 => x"d40c9353",
   869 => x"805287fc",
   870 => x"80c15199",
   871 => x"fd2d80c6",
   872 => x"94088b38",
   873 => x"81ff0bd4",
   874 => x"0c81539b",
   875 => x"b7049af0",
   876 => x"2dff1353",
   877 => x"72de3872",
   878 => x"80c6940c",
   879 => x"028c050d",
   880 => x"0402ec05",
   881 => x"0d810b80",
   882 => x"c6f80c84",
   883 => x"54d00870",
   884 => x"8f2a7081",
   885 => x"06515153",
   886 => x"72f33872",
   887 => x"d00c9af0",
   888 => x"2dbdc851",
   889 => x"86a02dd0",
   890 => x"08708f2a",
   891 => x"70810651",
   892 => x"515372f3",
   893 => x"38810bd0",
   894 => x"0cb15380",
   895 => x"5284d480",
   896 => x"c05199fd",
   897 => x"2d80c694",
   898 => x"08812e93",
   899 => x"3872822e",
   900 => x"bf38ff13",
   901 => x"5372e438",
   902 => x"ff145473",
   903 => x"ffaf389a",
   904 => x"f02d83aa",
   905 => x"52849c80",
   906 => x"c85199fd",
   907 => x"2d80c694",
   908 => x"08812e09",
   909 => x"81069338",
   910 => x"99ae2d80",
   911 => x"c6940883",
   912 => x"ffff0653",
   913 => x"7283aa2e",
   914 => x"9d389b89",
   915 => x"2d9ce104",
   916 => x"bdd45186",
   917 => x"a02d8053",
   918 => x"9eb604bd",
   919 => x"ec5186a0",
   920 => x"2d80549e",
   921 => x"870481ff",
   922 => x"0bd40cb1",
   923 => x"549af02d",
   924 => x"8fcf5380",
   925 => x"5287fc80",
   926 => x"f75199fd",
   927 => x"2d80c694",
   928 => x"085580c6",
   929 => x"9408812e",
   930 => x"0981069c",
   931 => x"3881ff0b",
   932 => x"d40c820a",
   933 => x"52849c80",
   934 => x"e95199fd",
   935 => x"2d80c694",
   936 => x"08802e8d",
   937 => x"389af02d",
   938 => x"ff135372",
   939 => x"c6389dfa",
   940 => x"0481ff0b",
   941 => x"d40c80c6",
   942 => x"94085287",
   943 => x"fc80fa51",
   944 => x"99fd2d80",
   945 => x"c69408b2",
   946 => x"3881ff0b",
   947 => x"d40cd408",
   948 => x"5381ff0b",
   949 => x"d40c81ff",
   950 => x"0bd40c81",
   951 => x"ff0bd40c",
   952 => x"81ff0bd4",
   953 => x"0c72862a",
   954 => x"70810676",
   955 => x"56515372",
   956 => x"963880c6",
   957 => x"9408549e",
   958 => x"87047382",
   959 => x"2efedc38",
   960 => x"ff145473",
   961 => x"fee73873",
   962 => x"80c6f80c",
   963 => x"738b3881",
   964 => x"5287fc80",
   965 => x"d05199fd",
   966 => x"2d81ff0b",
   967 => x"d40cd008",
   968 => x"708f2a70",
   969 => x"81065151",
   970 => x"5372f338",
   971 => x"72d00c81",
   972 => x"ff0bd40c",
   973 => x"81537280",
   974 => x"c6940c02",
   975 => x"94050d04",
   976 => x"02e8050d",
   977 => x"78558056",
   978 => x"81ff0bd4",
   979 => x"0cd00870",
   980 => x"8f2a7081",
   981 => x"06515153",
   982 => x"72f33882",
   983 => x"810bd00c",
   984 => x"81ff0bd4",
   985 => x"0c775287",
   986 => x"fc80d151",
   987 => x"99fd2d80",
   988 => x"dbc6df54",
   989 => x"80c69408",
   990 => x"802e8a38",
   991 => x"be8c5186",
   992 => x"a02d9fd9",
   993 => x"0481ff0b",
   994 => x"d40cd408",
   995 => x"7081ff06",
   996 => x"51537281",
   997 => x"fe2e0981",
   998 => x"069e3880",
   999 => x"ff5399ae",
  1000 => x"2d80c694",
  1001 => x"08757084",
  1002 => x"05570cff",
  1003 => x"13537280",
  1004 => x"25ec3881",
  1005 => x"569fbe04",
  1006 => x"ff145473",
  1007 => x"c83881ff",
  1008 => x"0bd40c81",
  1009 => x"ff0bd40c",
  1010 => x"d008708f",
  1011 => x"2a708106",
  1012 => x"51515372",
  1013 => x"f33872d0",
  1014 => x"0c7580c6",
  1015 => x"940c0298",
  1016 => x"050d0402",
  1017 => x"e8050d77",
  1018 => x"797b5855",
  1019 => x"55805372",
  1020 => x"7625a338",
  1021 => x"74708105",
  1022 => x"5680f52d",
  1023 => x"74708105",
  1024 => x"5680f52d",
  1025 => x"52527171",
  1026 => x"2e863881",
  1027 => x"51a09804",
  1028 => x"8113539f",
  1029 => x"ef048051",
  1030 => x"7080c694",
  1031 => x"0c029805",
  1032 => x"0d0402ec",
  1033 => x"050d7655",
  1034 => x"74802e80",
  1035 => x"c2389a15",
  1036 => x"80e02d51",
  1037 => x"aeaf2d80",
  1038 => x"c6940880",
  1039 => x"c6940880",
  1040 => x"cdac0c80",
  1041 => x"c6940854",
  1042 => x"5480cd88",
  1043 => x"08802e9a",
  1044 => x"38941580",
  1045 => x"e02d51ae",
  1046 => x"af2d80c6",
  1047 => x"9408902b",
  1048 => x"83fff00a",
  1049 => x"06707507",
  1050 => x"51537280",
  1051 => x"cdac0c80",
  1052 => x"cdac0853",
  1053 => x"72802e9d",
  1054 => x"3880cd80",
  1055 => x"08fe1471",
  1056 => x"2980cd94",
  1057 => x"080580cd",
  1058 => x"b00c7084",
  1059 => x"2b80cd8c",
  1060 => x"0c54a1c3",
  1061 => x"0480cd98",
  1062 => x"0880cdac",
  1063 => x"0c80cd9c",
  1064 => x"0880cdb0",
  1065 => x"0c80cd88",
  1066 => x"08802e8b",
  1067 => x"3880cd80",
  1068 => x"08842b53",
  1069 => x"a1be0480",
  1070 => x"cda00884",
  1071 => x"2b537280",
  1072 => x"cd8c0c02",
  1073 => x"94050d04",
  1074 => x"02d8050d",
  1075 => x"800b80cd",
  1076 => x"880c8454",
  1077 => x"9bc12d80",
  1078 => x"c6940880",
  1079 => x"2e973880",
  1080 => x"c6fc5280",
  1081 => x"519ec02d",
  1082 => x"80c69408",
  1083 => x"802e8638",
  1084 => x"fe54a1fd",
  1085 => x"04ff1454",
  1086 => x"738024d8",
  1087 => x"38738c38",
  1088 => x"be9c5186",
  1089 => x"a02d7355",
  1090 => x"a7ca0480",
  1091 => x"56810b80",
  1092 => x"cdb40c88",
  1093 => x"53beb052",
  1094 => x"80c7b251",
  1095 => x"9fe32d80",
  1096 => x"c6940876",
  1097 => x"2e098106",
  1098 => x"893880c6",
  1099 => x"940880cd",
  1100 => x"b40c8853",
  1101 => x"bebc5280",
  1102 => x"c7ce519f",
  1103 => x"e32d80c6",
  1104 => x"94088938",
  1105 => x"80c69408",
  1106 => x"80cdb40c",
  1107 => x"80cdb408",
  1108 => x"802e8180",
  1109 => x"3880cac2",
  1110 => x"0b80f52d",
  1111 => x"80cac30b",
  1112 => x"80f52d71",
  1113 => x"982b7190",
  1114 => x"2b0780ca",
  1115 => x"c40b80f5",
  1116 => x"2d70882b",
  1117 => x"720780ca",
  1118 => x"c50b80f5",
  1119 => x"2d710780",
  1120 => x"cafa0b80",
  1121 => x"f52d80ca",
  1122 => x"fb0b80f5",
  1123 => x"2d71882b",
  1124 => x"07535f54",
  1125 => x"525a5657",
  1126 => x"557381ab",
  1127 => x"aa2e0981",
  1128 => x"068e3875",
  1129 => x"51adfe2d",
  1130 => x"80c69408",
  1131 => x"56a3bd04",
  1132 => x"7382d4d5",
  1133 => x"2e8738be",
  1134 => x"c851a486",
  1135 => x"0480c6fc",
  1136 => x"5275519e",
  1137 => x"c02d80c6",
  1138 => x"94085580",
  1139 => x"c6940880",
  1140 => x"2e83f738",
  1141 => x"8853bebc",
  1142 => x"5280c7ce",
  1143 => x"519fe32d",
  1144 => x"80c69408",
  1145 => x"8a38810b",
  1146 => x"80cd880c",
  1147 => x"a48c0488",
  1148 => x"53beb052",
  1149 => x"80c7b251",
  1150 => x"9fe32d80",
  1151 => x"c6940880",
  1152 => x"2e8a38be",
  1153 => x"dc5186a0",
  1154 => x"2da4eb04",
  1155 => x"80cafa0b",
  1156 => x"80f52d54",
  1157 => x"7380d52e",
  1158 => x"09810680",
  1159 => x"ce3880ca",
  1160 => x"fb0b80f5",
  1161 => x"2d547381",
  1162 => x"aa2e0981",
  1163 => x"06bd3880",
  1164 => x"0b80c6fc",
  1165 => x"0b80f52d",
  1166 => x"56547481",
  1167 => x"e92e8338",
  1168 => x"81547481",
  1169 => x"eb2e8c38",
  1170 => x"80557375",
  1171 => x"2e098106",
  1172 => x"82f83880",
  1173 => x"c7870b80",
  1174 => x"f52d5574",
  1175 => x"8e3880c7",
  1176 => x"880b80f5",
  1177 => x"2d547382",
  1178 => x"2e863880",
  1179 => x"55a7ca04",
  1180 => x"80c7890b",
  1181 => x"80f52d70",
  1182 => x"80cd800c",
  1183 => x"ff0580cd",
  1184 => x"840c80c7",
  1185 => x"8a0b80f5",
  1186 => x"2d80c78b",
  1187 => x"0b80f52d",
  1188 => x"58760577",
  1189 => x"82802905",
  1190 => x"7080cd90",
  1191 => x"0c80c78c",
  1192 => x"0b80f52d",
  1193 => x"7080cda4",
  1194 => x"0c80cd88",
  1195 => x"08595758",
  1196 => x"76802e81",
  1197 => x"b6388853",
  1198 => x"bebc5280",
  1199 => x"c7ce519f",
  1200 => x"e32d80c6",
  1201 => x"94088282",
  1202 => x"3880cd80",
  1203 => x"0870842b",
  1204 => x"80cd8c0c",
  1205 => x"7080cda0",
  1206 => x"0c80c7a1",
  1207 => x"0b80f52d",
  1208 => x"80c7a00b",
  1209 => x"80f52d71",
  1210 => x"82802905",
  1211 => x"80c7a20b",
  1212 => x"80f52d70",
  1213 => x"84808029",
  1214 => x"1280c7a3",
  1215 => x"0b80f52d",
  1216 => x"7081800a",
  1217 => x"29127080",
  1218 => x"cda80c80",
  1219 => x"cda40871",
  1220 => x"2980cd90",
  1221 => x"08057080",
  1222 => x"cd940c80",
  1223 => x"c7a90b80",
  1224 => x"f52d80c7",
  1225 => x"a80b80f5",
  1226 => x"2d718280",
  1227 => x"290580c7",
  1228 => x"aa0b80f5",
  1229 => x"2d708480",
  1230 => x"80291280",
  1231 => x"c7ab0b80",
  1232 => x"f52d7098",
  1233 => x"2b81f00a",
  1234 => x"06720570",
  1235 => x"80cd980c",
  1236 => x"fe117e29",
  1237 => x"770580cd",
  1238 => x"9c0c5259",
  1239 => x"5243545e",
  1240 => x"51525952",
  1241 => x"5d575957",
  1242 => x"a7c30480",
  1243 => x"c78e0b80",
  1244 => x"f52d80c7",
  1245 => x"8d0b80f5",
  1246 => x"2d718280",
  1247 => x"29057080",
  1248 => x"cd8c0c70",
  1249 => x"a02983ff",
  1250 => x"0570892a",
  1251 => x"7080cda0",
  1252 => x"0c80c793",
  1253 => x"0b80f52d",
  1254 => x"80c7920b",
  1255 => x"80f52d71",
  1256 => x"82802905",
  1257 => x"7080cda8",
  1258 => x"0c7b7129",
  1259 => x"1e7080cd",
  1260 => x"9c0c7d80",
  1261 => x"cd980c73",
  1262 => x"0580cd94",
  1263 => x"0c555e51",
  1264 => x"51555580",
  1265 => x"51a0a22d",
  1266 => x"81557480",
  1267 => x"c6940c02",
  1268 => x"a8050d04",
  1269 => x"02ec050d",
  1270 => x"7670872c",
  1271 => x"7180ff06",
  1272 => x"55565480",
  1273 => x"cd88088a",
  1274 => x"3873882c",
  1275 => x"7481ff06",
  1276 => x"545580c6",
  1277 => x"fc5280cd",
  1278 => x"90081551",
  1279 => x"9ec02d80",
  1280 => x"c6940854",
  1281 => x"80c69408",
  1282 => x"802eb838",
  1283 => x"80cd8808",
  1284 => x"802e9a38",
  1285 => x"72842980",
  1286 => x"c6fc0570",
  1287 => x"085253ad",
  1288 => x"fe2d80c6",
  1289 => x"9408f00a",
  1290 => x"0653a8c1",
  1291 => x"04721080",
  1292 => x"c6fc0570",
  1293 => x"80e02d52",
  1294 => x"53aeaf2d",
  1295 => x"80c69408",
  1296 => x"53725473",
  1297 => x"80c6940c",
  1298 => x"0294050d",
  1299 => x"0402e005",
  1300 => x"0d797084",
  1301 => x"2c80cdb0",
  1302 => x"0805718f",
  1303 => x"06525553",
  1304 => x"728a3880",
  1305 => x"c6fc5273",
  1306 => x"519ec02d",
  1307 => x"72a02980",
  1308 => x"c6fc0554",
  1309 => x"807480f5",
  1310 => x"2d565374",
  1311 => x"732e8338",
  1312 => x"81537481",
  1313 => x"e52e81f4",
  1314 => x"38817074",
  1315 => x"06545872",
  1316 => x"802e81e8",
  1317 => x"388b1480",
  1318 => x"f52d7083",
  1319 => x"2a790658",
  1320 => x"56769b38",
  1321 => x"80c4d808",
  1322 => x"53728938",
  1323 => x"7280cafc",
  1324 => x"0b81b72d",
  1325 => x"7680c4d8",
  1326 => x"0c7353aa",
  1327 => x"fe04758f",
  1328 => x"2e098106",
  1329 => x"81b63874",
  1330 => x"9f068d29",
  1331 => x"80caef11",
  1332 => x"51538114",
  1333 => x"80f52d73",
  1334 => x"70810555",
  1335 => x"81b72d83",
  1336 => x"1480f52d",
  1337 => x"73708105",
  1338 => x"5581b72d",
  1339 => x"851480f5",
  1340 => x"2d737081",
  1341 => x"055581b7",
  1342 => x"2d871480",
  1343 => x"f52d7370",
  1344 => x"81055581",
  1345 => x"b72d8914",
  1346 => x"80f52d73",
  1347 => x"70810555",
  1348 => x"81b72d8e",
  1349 => x"1480f52d",
  1350 => x"73708105",
  1351 => x"5581b72d",
  1352 => x"901480f5",
  1353 => x"2d737081",
  1354 => x"055581b7",
  1355 => x"2d921480",
  1356 => x"f52d7370",
  1357 => x"81055581",
  1358 => x"b72d9414",
  1359 => x"80f52d73",
  1360 => x"70810555",
  1361 => x"81b72d96",
  1362 => x"1480f52d",
  1363 => x"73708105",
  1364 => x"5581b72d",
  1365 => x"981480f5",
  1366 => x"2d737081",
  1367 => x"055581b7",
  1368 => x"2d9c1480",
  1369 => x"f52d7370",
  1370 => x"81055581",
  1371 => x"b72d9e14",
  1372 => x"80f52d73",
  1373 => x"81b72d77",
  1374 => x"80c4d80c",
  1375 => x"80537280",
  1376 => x"c6940c02",
  1377 => x"a0050d04",
  1378 => x"02cc050d",
  1379 => x"7e605e5a",
  1380 => x"800b80cd",
  1381 => x"ac0880cd",
  1382 => x"b008595c",
  1383 => x"56805880",
  1384 => x"cd8c0878",
  1385 => x"2e81b838",
  1386 => x"778f06a0",
  1387 => x"17575473",
  1388 => x"913880c6",
  1389 => x"fc527651",
  1390 => x"8117579e",
  1391 => x"c02d80c6",
  1392 => x"fc568076",
  1393 => x"80f52d56",
  1394 => x"5474742e",
  1395 => x"83388154",
  1396 => x"7481e52e",
  1397 => x"80fd3881",
  1398 => x"70750655",
  1399 => x"5c73802e",
  1400 => x"80f1388b",
  1401 => x"1680f52d",
  1402 => x"98065978",
  1403 => x"80e5388b",
  1404 => x"537c5275",
  1405 => x"519fe32d",
  1406 => x"80c69408",
  1407 => x"80d5389c",
  1408 => x"160851ad",
  1409 => x"fe2d80c6",
  1410 => x"9408841b",
  1411 => x"0c9a1680",
  1412 => x"e02d51ae",
  1413 => x"af2d80c6",
  1414 => x"940880c6",
  1415 => x"9408881c",
  1416 => x"0c80c694",
  1417 => x"08555580",
  1418 => x"cd880880",
  1419 => x"2e993894",
  1420 => x"1680e02d",
  1421 => x"51aeaf2d",
  1422 => x"80c69408",
  1423 => x"902b83ff",
  1424 => x"f00a0670",
  1425 => x"16515473",
  1426 => x"881b0c78",
  1427 => x"7a0c7b54",
  1428 => x"ad9b0481",
  1429 => x"185880cd",
  1430 => x"8c087826",
  1431 => x"feca3880",
  1432 => x"cd880880",
  1433 => x"2eb3387a",
  1434 => x"51a7d42d",
  1435 => x"80c69408",
  1436 => x"80c69408",
  1437 => x"80ffffff",
  1438 => x"f806555b",
  1439 => x"7380ffff",
  1440 => x"fff82e95",
  1441 => x"3880c694",
  1442 => x"08fe0580",
  1443 => x"cd800829",
  1444 => x"80cd9408",
  1445 => x"0557ab9d",
  1446 => x"04805473",
  1447 => x"80c6940c",
  1448 => x"02b4050d",
  1449 => x"0402f405",
  1450 => x"0d747008",
  1451 => x"8105710c",
  1452 => x"700880cd",
  1453 => x"84080653",
  1454 => x"53718f38",
  1455 => x"88130851",
  1456 => x"a7d42d80",
  1457 => x"c6940888",
  1458 => x"140c810b",
  1459 => x"80c6940c",
  1460 => x"028c050d",
  1461 => x"0402f005",
  1462 => x"0d758811",
  1463 => x"08fe0580",
  1464 => x"cd800829",
  1465 => x"80cd9408",
  1466 => x"11720880",
  1467 => x"cd840806",
  1468 => x"05795553",
  1469 => x"54549ec0",
  1470 => x"2d029005",
  1471 => x"0d0402f4",
  1472 => x"050d7470",
  1473 => x"882a83fe",
  1474 => x"80067072",
  1475 => x"982a0772",
  1476 => x"882b87fc",
  1477 => x"80800673",
  1478 => x"982b81f0",
  1479 => x"0a067173",
  1480 => x"070780c6",
  1481 => x"940c5651",
  1482 => x"5351028c",
  1483 => x"050d0402",
  1484 => x"f8050d02",
  1485 => x"8e0580f5",
  1486 => x"2d74882b",
  1487 => x"077083ff",
  1488 => x"ff0680c6",
  1489 => x"940c5102",
  1490 => x"88050d04",
  1491 => x"02f4050d",
  1492 => x"74767853",
  1493 => x"54528071",
  1494 => x"25973872",
  1495 => x"70810554",
  1496 => x"80f52d72",
  1497 => x"70810554",
  1498 => x"81b72dff",
  1499 => x"115170eb",
  1500 => x"38807281",
  1501 => x"b72d028c",
  1502 => x"050d0402",
  1503 => x"e8050d77",
  1504 => x"56807056",
  1505 => x"54737624",
  1506 => x"b63880cd",
  1507 => x"8c08742e",
  1508 => x"ae387351",
  1509 => x"a8cd2d80",
  1510 => x"c6940880",
  1511 => x"c6940809",
  1512 => x"81057080",
  1513 => x"c6940807",
  1514 => x"9f2a7705",
  1515 => x"81175757",
  1516 => x"53537476",
  1517 => x"24893880",
  1518 => x"cd8c0874",
  1519 => x"26d43872",
  1520 => x"80c6940c",
  1521 => x"0298050d",
  1522 => x"0402f005",
  1523 => x"0d80c690",
  1524 => x"081651ae",
  1525 => x"fb2d80c6",
  1526 => x"9408802e",
  1527 => x"9f388b53",
  1528 => x"80c69408",
  1529 => x"5280cafc",
  1530 => x"51aecc2d",
  1531 => x"80cdb808",
  1532 => x"5473802e",
  1533 => x"873880ca",
  1534 => x"fc51732d",
  1535 => x"0290050d",
  1536 => x"0402dc05",
  1537 => x"0d80705a",
  1538 => x"557480c6",
  1539 => x"900825b4",
  1540 => x"3880cd8c",
  1541 => x"08752eac",
  1542 => x"387851a8",
  1543 => x"cd2d80c6",
  1544 => x"94080981",
  1545 => x"057080c6",
  1546 => x"9408079f",
  1547 => x"2a760581",
  1548 => x"1b5b5654",
  1549 => x"7480c690",
  1550 => x"08258938",
  1551 => x"80cd8c08",
  1552 => x"7926d638",
  1553 => x"80557880",
  1554 => x"cd8c0827",
  1555 => x"81db3878",
  1556 => x"51a8cd2d",
  1557 => x"80c69408",
  1558 => x"802e81ad",
  1559 => x"3880c694",
  1560 => x"088b0580",
  1561 => x"f52d7084",
  1562 => x"2a708106",
  1563 => x"77107884",
  1564 => x"2b80cafc",
  1565 => x"0b80f52d",
  1566 => x"5c5c5351",
  1567 => x"55567380",
  1568 => x"2e80cb38",
  1569 => x"7416822b",
  1570 => x"b2cd0b80",
  1571 => x"c4e4120c",
  1572 => x"54777531",
  1573 => x"1080cdbc",
  1574 => x"11555690",
  1575 => x"74708105",
  1576 => x"5681b72d",
  1577 => x"a07481b7",
  1578 => x"2d7681ff",
  1579 => x"06811658",
  1580 => x"5473802e",
  1581 => x"8a389c53",
  1582 => x"80cafc52",
  1583 => x"b1c6048b",
  1584 => x"5380c694",
  1585 => x"085280cd",
  1586 => x"be1651b2",
  1587 => x"81047416",
  1588 => x"822bafc9",
  1589 => x"0b80c4e4",
  1590 => x"120c5476",
  1591 => x"81ff0681",
  1592 => x"16585473",
  1593 => x"802e8a38",
  1594 => x"9c5380ca",
  1595 => x"fc52b1f8",
  1596 => x"048b5380",
  1597 => x"c6940852",
  1598 => x"77753110",
  1599 => x"80cdbc05",
  1600 => x"517655ae",
  1601 => x"cc2db29e",
  1602 => x"04749029",
  1603 => x"75317010",
  1604 => x"80cdbc05",
  1605 => x"515480c6",
  1606 => x"94087481",
  1607 => x"b72d8119",
  1608 => x"59748b24",
  1609 => x"a338b0c6",
  1610 => x"04749029",
  1611 => x"75317010",
  1612 => x"80cdbc05",
  1613 => x"8c773157",
  1614 => x"51548074",
  1615 => x"81b72d9e",
  1616 => x"14ff1656",
  1617 => x"5474f338",
  1618 => x"02a4050d",
  1619 => x"0402fc05",
  1620 => x"0d80c690",
  1621 => x"081351ae",
  1622 => x"fb2d80c6",
  1623 => x"9408802e",
  1624 => x"893880c6",
  1625 => x"940851a0",
  1626 => x"a22d800b",
  1627 => x"80c6900c",
  1628 => x"b0812d91",
  1629 => x"892d0284",
  1630 => x"050d0402",
  1631 => x"fc050d72",
  1632 => x"5170fd2e",
  1633 => x"b03870fd",
  1634 => x"248a3870",
  1635 => x"fc2e80cc",
  1636 => x"38b3e604",
  1637 => x"70fe2eb7",
  1638 => x"3870ff2e",
  1639 => x"09810680",
  1640 => x"c53880c6",
  1641 => x"90085170",
  1642 => x"802ebb38",
  1643 => x"ff1180c6",
  1644 => x"900cb3e6",
  1645 => x"0480c690",
  1646 => x"08f00570",
  1647 => x"80c6900c",
  1648 => x"51708025",
  1649 => x"a138800b",
  1650 => x"80c6900c",
  1651 => x"b3e60480",
  1652 => x"c6900881",
  1653 => x"0580c690",
  1654 => x"0cb3e604",
  1655 => x"80c69008",
  1656 => x"900580c6",
  1657 => x"900cb081",
  1658 => x"2d91892d",
  1659 => x"0284050d",
  1660 => x"0402fc05",
  1661 => x"0d800b80",
  1662 => x"c6900cb0",
  1663 => x"812d9099",
  1664 => x"2d80c694",
  1665 => x"0880c680",
  1666 => x"0c80c4dc",
  1667 => x"5192ac2d",
  1668 => x"0284050d",
  1669 => x"047180cd",
  1670 => x"b80c0400",
  1671 => x"00ffffff",
  1672 => x"ff00ffff",
  1673 => x"ffff00ff",
  1674 => x"ffffff00",
  1675 => x"45786974",
  1676 => x"00000000",
  1677 => x"506f7420",
  1678 => x"33263420",
  1679 => x"4a6f7920",
  1680 => x"32204469",
  1681 => x"73706172",
  1682 => x"6f20322f",
  1683 => x"33000000",
  1684 => x"506f7420",
  1685 => x"33263420",
  1686 => x"5261746f",
  1687 => x"6e000000",
  1688 => x"506f7420",
  1689 => x"33263420",
  1690 => x"50616464",
  1691 => x"6c657320",
  1692 => x"33263400",
  1693 => x"506f7420",
  1694 => x"31263220",
  1695 => x"4a6f7920",
  1696 => x"31204469",
  1697 => x"73706172",
  1698 => x"6f20322f",
  1699 => x"33000000",
  1700 => x"506f7420",
  1701 => x"31263220",
  1702 => x"5261746f",
  1703 => x"6e000000",
  1704 => x"506f7420",
  1705 => x"31263220",
  1706 => x"50616464",
  1707 => x"6c657320",
  1708 => x"31263200",
  1709 => x"50756572",
  1710 => x"746f2055",
  1711 => x"41525400",
  1712 => x"50756572",
  1713 => x"746f204a",
  1714 => x"6f797374",
  1715 => x"69636b73",
  1716 => x"00000000",
  1717 => x"4a6f7973",
  1718 => x"7469636b",
  1719 => x"73204e6f",
  1720 => x"726d616c",
  1721 => x"00000000",
  1722 => x"4a6f7973",
  1723 => x"7469636b",
  1724 => x"7320496e",
  1725 => x"74657263",
  1726 => x"616d6269",
  1727 => x"61646f73",
  1728 => x"00000000",
  1729 => x"4d657a63",
  1730 => x"6c612053",
  1731 => x"74657265",
  1732 => x"6f204e6f",
  1733 => x"00000000",
  1734 => x"4d657a63",
  1735 => x"6c612053",
  1736 => x"74657265",
  1737 => x"6f203235",
  1738 => x"25000000",
  1739 => x"4d657a63",
  1740 => x"6c612053",
  1741 => x"74657265",
  1742 => x"6f203530",
  1743 => x"25000000",
  1744 => x"4d657a63",
  1745 => x"6c612053",
  1746 => x"74657265",
  1747 => x"6f203735",
  1748 => x"25000000",
  1749 => x"45787061",
  1750 => x"6e73696f",
  1751 => x"6e206465",
  1752 => x"20536f6e",
  1753 => x"69646f20",
  1754 => x"4e6f0000",
  1755 => x"45787061",
  1756 => x"6e73696f",
  1757 => x"6e206465",
  1758 => x"20536f6e",
  1759 => x"69646f20",
  1760 => x"4f504c32",
  1761 => x"00000000",
  1762 => x"46696c74",
  1763 => x"726f2064",
  1764 => x"65204175",
  1765 => x"64696f20",
  1766 => x"4f6e0000",
  1767 => x"46696c74",
  1768 => x"726f2064",
  1769 => x"65204175",
  1770 => x"64696f20",
  1771 => x"4f666600",
  1772 => x"53494420",
  1773 => x"44657265",
  1774 => x"63686f20",
  1775 => x"41646472",
  1776 => x"20496775",
  1777 => x"616c0000",
  1778 => x"53494420",
  1779 => x"44657265",
  1780 => x"63686f20",
  1781 => x"41646472",
  1782 => x"20444530",
  1783 => x"30000000",
  1784 => x"53494420",
  1785 => x"44657265",
  1786 => x"63686f20",
  1787 => x"41646472",
  1788 => x"20443432",
  1789 => x"30000000",
  1790 => x"53494420",
  1791 => x"44657265",
  1792 => x"63686f20",
  1793 => x"41646472",
  1794 => x"20443530",
  1795 => x"30000000",
  1796 => x"53494420",
  1797 => x"44657265",
  1798 => x"63686f20",
  1799 => x"41646472",
  1800 => x"20444630",
  1801 => x"30000000",
  1802 => x"53494420",
  1803 => x"44657265",
  1804 => x"63686f20",
  1805 => x"36353831",
  1806 => x"00000000",
  1807 => x"53494420",
  1808 => x"44657265",
  1809 => x"63686f20",
  1810 => x"38353830",
  1811 => x"00000000",
  1812 => x"53494420",
  1813 => x"497a7175",
  1814 => x"69657264",
  1815 => x"6f203635",
  1816 => x"38310000",
  1817 => x"53494420",
  1818 => x"497a7175",
  1819 => x"69657264",
  1820 => x"6f203835",
  1821 => x"38300000",
  1822 => x"5363616e",
  1823 => x"646f7562",
  1824 => x"6c657220",
  1825 => x"4e696e67",
  1826 => x"756e6f00",
  1827 => x"5363616e",
  1828 => x"646f7562",
  1829 => x"6c657220",
  1830 => x"48513278",
  1831 => x"2d333230",
  1832 => x"00000000",
  1833 => x"5363616e",
  1834 => x"646f7562",
  1835 => x"6c657220",
  1836 => x"48513278",
  1837 => x"2d313630",
  1838 => x"00000000",
  1839 => x"5363616e",
  1840 => x"646f7562",
  1841 => x"6c657220",
  1842 => x"43525420",
  1843 => x"32352500",
  1844 => x"5363616e",
  1845 => x"646f7562",
  1846 => x"6c657220",
  1847 => x"43525420",
  1848 => x"35302500",
  1849 => x"5363616e",
  1850 => x"646f7562",
  1851 => x"6c657220",
  1852 => x"43525420",
  1853 => x"37352500",
  1854 => x"466f726d",
  1855 => x"61746f20",
  1856 => x"4f726967",
  1857 => x"696e616c",
  1858 => x"00000000",
  1859 => x"466f726d",
  1860 => x"61746f20",
  1861 => x"50616e74",
  1862 => x"616c6c61",
  1863 => x"20436f6d",
  1864 => x"706c6574",
  1865 => x"61000000",
  1866 => x"466f726d",
  1867 => x"61746f20",
  1868 => x"5b415243",
  1869 => x"315d0000",
  1870 => x"466f726d",
  1871 => x"61746f20",
  1872 => x"5b415243",
  1873 => x"325d0000",
  1874 => x"41737065",
  1875 => x"63746f20",
  1876 => x"4f726967",
  1877 => x"696e616c",
  1878 => x"00000000",
  1879 => x"41737065",
  1880 => x"63746f20",
  1881 => x"416e6368",
  1882 => x"6f000000",
  1883 => x"56696465",
  1884 => x"6f205041",
  1885 => x"4c000000",
  1886 => x"56696465",
  1887 => x"6f204e54",
  1888 => x"53430000",
  1889 => x"2020203d",
  1890 => x"434f4d4f",
  1891 => x"444f5245",
  1892 => x"2036343d",
  1893 => x"20202000",
  1894 => x"20202062",
  1895 => x"79204e65",
  1896 => x"75726f52",
  1897 => x"756c657a",
  1898 => x"20202000",
  1899 => x"20202020",
  1900 => x"20202020",
  1901 => x"20202020",
  1902 => x"20202020",
  1903 => x"20202000",
  1904 => x"52657365",
  1905 => x"74000000",
  1906 => x"52657365",
  1907 => x"74202620",
  1908 => x"536f6c74",
  1909 => x"61722043",
  1910 => x"61727475",
  1911 => x"63686f00",
  1912 => x"56696465",
  1913 => x"6f201000",
  1914 => x"41756469",
  1915 => x"6f201000",
  1916 => x"50756572",
  1917 => x"746f7320",
  1918 => x"10000000",
  1919 => x"53616361",
  1920 => x"72204369",
  1921 => x"6e746100",
  1922 => x"506c6179",
  1923 => x"2f53746f",
  1924 => x"70204369",
  1925 => x"6e746100",
  1926 => x"43617267",
  1927 => x"61722044",
  1928 => x"6973636f",
  1929 => x"2f43696e",
  1930 => x"74612f43",
  1931 => x"61727420",
  1932 => x"10000000",
  1933 => x"44697363",
  1934 => x"6f204772",
  1935 => x"61626162",
  1936 => x"6c650000",
  1937 => x"44697363",
  1938 => x"6f20536f",
  1939 => x"6c6f204c",
  1940 => x"65637475",
  1941 => x"72610000",
  1942 => x"536f6e69",
  1943 => x"646f2043",
  1944 => x"696e7461",
  1945 => x"204f6666",
  1946 => x"00000000",
  1947 => x"536f6e69",
  1948 => x"646f2043",
  1949 => x"696e7461",
  1950 => x"204f6e00",
  1951 => x"4b65726e",
  1952 => x"656c2043",
  1953 => x"61726761",
  1954 => x"626c6500",
  1955 => x"4b65726e",
  1956 => x"656c2043",
  1957 => x"36340000",
  1958 => x"4b65726e",
  1959 => x"656c2043",
  1960 => x"36344753",
  1961 => x"00000000",
  1962 => x"43617267",
  1963 => x"61204661",
  1964 => x"6c6c6964",
  1965 => x"61000000",
  1966 => x"4f4b0000",
  1967 => x"16200000",
  1968 => x"14200000",
  1969 => x"15200000",
  1970 => x"53442069",
  1971 => x"6e69742e",
  1972 => x"2e2e0a00",
  1973 => x"53442063",
  1974 => x"61726420",
  1975 => x"72657365",
  1976 => x"74206661",
  1977 => x"696c6564",
  1978 => x"210a0000",
  1979 => x"53444843",
  1980 => x"20657272",
  1981 => x"6f72210a",
  1982 => x"00000000",
  1983 => x"57726974",
  1984 => x"65206661",
  1985 => x"696c6564",
  1986 => x"0a000000",
  1987 => x"52656164",
  1988 => x"20666169",
  1989 => x"6c65640a",
  1990 => x"00000000",
  1991 => x"43617264",
  1992 => x"20696e69",
  1993 => x"74206661",
  1994 => x"696c6564",
  1995 => x"0a000000",
  1996 => x"46415431",
  1997 => x"36202020",
  1998 => x"00000000",
  1999 => x"46415433",
  2000 => x"32202020",
  2001 => x"00000000",
  2002 => x"4e6f2070",
  2003 => x"61727469",
  2004 => x"74696f6e",
  2005 => x"20736967",
  2006 => x"0a000000",
  2007 => x"42616420",
  2008 => x"70617274",
  2009 => x"0a000000",
  2010 => x"4261636b",
  2011 => x"00000000",
  2012 => x"00000002",
  2013 => x"00000003",
  2014 => x"00001fdc",
  2015 => x"00000002",
  2016 => x"00000003",
  2017 => x"00001fd4",
  2018 => x"00000002",
  2019 => x"00000003",
  2020 => x"00001fc8",
  2021 => x"00000003",
  2022 => x"00000003",
  2023 => x"00001fbc",
  2024 => x"00000003",
  2025 => x"00000004",
  2026 => x"00001a2c",
  2027 => x"00002108",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00000000",
  2031 => x"00001a34",
  2032 => x"00001a50",
  2033 => x"00001a60",
  2034 => x"00001a74",
  2035 => x"00001a90",
  2036 => x"00001aa0",
  2037 => x"00001ab4",
  2038 => x"00001ac0",
  2039 => x"00001ad4",
  2040 => x"00001ae8",
  2041 => x"00000003",
  2042 => x"00002080",
  2043 => x"00000002",
  2044 => x"00000003",
  2045 => x"00002078",
  2046 => x"00000002",
  2047 => x"00000003",
  2048 => x"00002064",
  2049 => x"00000005",
  2050 => x"00000003",
  2051 => x"0000205c",
  2052 => x"00000002",
  2053 => x"00000003",
  2054 => x"00002054",
  2055 => x"00000002",
  2056 => x"00000003",
  2057 => x"00002044",
  2058 => x"00000004",
  2059 => x"00000004",
  2060 => x"00001a2c",
  2061 => x"00002108",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00001b04",
  2066 => x"00001b18",
  2067 => x"00001b2c",
  2068 => x"00001b40",
  2069 => x"00001b54",
  2070 => x"00001b6c",
  2071 => x"00001b88",
  2072 => x"00001b9c",
  2073 => x"00001bb0",
  2074 => x"00001bc8",
  2075 => x"00001be0",
  2076 => x"00001bf8",
  2077 => x"00001c10",
  2078 => x"00001c28",
  2079 => x"00001c3c",
  2080 => x"00001c50",
  2081 => x"00001c64",
  2082 => x"00000003",
  2083 => x"00002100",
  2084 => x"00000002",
  2085 => x"00000003",
  2086 => x"000020f8",
  2087 => x"00000002",
  2088 => x"00000003",
  2089 => x"000020e8",
  2090 => x"00000004",
  2091 => x"00000003",
  2092 => x"000020d0",
  2093 => x"00000006",
  2094 => x"00000004",
  2095 => x"00001a2c",
  2096 => x"00002108",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00001c78",
  2101 => x"00001c8c",
  2102 => x"00001ca4",
  2103 => x"00001cbc",
  2104 => x"00001cd0",
  2105 => x"00001ce4",
  2106 => x"00001cf8",
  2107 => x"00001d0c",
  2108 => x"00001d28",
  2109 => x"00001d38",
  2110 => x"00001d48",
  2111 => x"00001d5c",
  2112 => x"00001d6c",
  2113 => x"00001d78",
  2114 => x"00000002",
  2115 => x"00001d84",
  2116 => x"00000000",
  2117 => x"00000002",
  2118 => x"00001d98",
  2119 => x"00000000",
  2120 => x"00000002",
  2121 => x"00001dac",
  2122 => x"00000000",
  2123 => x"00000002",
  2124 => x"00001dc0",
  2125 => x"00000371",
  2126 => x"00000002",
  2127 => x"00001dc8",
  2128 => x"00000388",
  2129 => x"00000004",
  2130 => x"00001de0",
  2131 => x"00002088",
  2132 => x"00000004",
  2133 => x"00001de8",
  2134 => x"00001fe4",
  2135 => x"00000004",
  2136 => x"00001df0",
  2137 => x"00001f74",
  2138 => x"00000003",
  2139 => x"000021d8",
  2140 => x"00000003",
  2141 => x"00000003",
  2142 => x"000021d0",
  2143 => x"00000002",
  2144 => x"00000003",
  2145 => x"000021c8",
  2146 => x"00000002",
  2147 => x"00000002",
  2148 => x"00001dfc",
  2149 => x"000003b8",
  2150 => x"00000002",
  2151 => x"00001e08",
  2152 => x"000003a0",
  2153 => x"00000002",
  2154 => x"00001e18",
  2155 => x"000019f1",
  2156 => x"00000002",
  2157 => x"00001a2c",
  2158 => x"00000822",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00001e34",
  2163 => x"00001e44",
  2164 => x"00001e58",
  2165 => x"00001e6c",
  2166 => x"00001e7c",
  2167 => x"00001e8c",
  2168 => x"00001e98",
  2169 => x"00000004",
  2170 => x"00001ea8",
  2171 => x"000021e4",
  2172 => x"00000004",
  2173 => x"00001eb8",
  2174 => x"00002108",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000002",
  2200 => x"000026bc",
  2201 => x"000017c9",
  2202 => x"00000002",
  2203 => x"000026da",
  2204 => x"000017c9",
  2205 => x"00000002",
  2206 => x"000026f8",
  2207 => x"000017c9",
  2208 => x"00000002",
  2209 => x"00002716",
  2210 => x"000017c9",
  2211 => x"00000002",
  2212 => x"00002734",
  2213 => x"000017c9",
  2214 => x"00000002",
  2215 => x"00002752",
  2216 => x"000017c9",
  2217 => x"00000002",
  2218 => x"00002770",
  2219 => x"000017c9",
  2220 => x"00000002",
  2221 => x"0000278e",
  2222 => x"000017c9",
  2223 => x"00000002",
  2224 => x"000027ac",
  2225 => x"000017c9",
  2226 => x"00000002",
  2227 => x"000027ca",
  2228 => x"000017c9",
  2229 => x"00000002",
  2230 => x"000027e8",
  2231 => x"000017c9",
  2232 => x"00000002",
  2233 => x"00002806",
  2234 => x"000017c9",
  2235 => x"00000002",
  2236 => x"00002824",
  2237 => x"000017c9",
  2238 => x"00000004",
  2239 => x"00001f68",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"0000197b",
  2244 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

