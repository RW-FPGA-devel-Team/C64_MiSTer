-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c7",
     9 => x"c4080b0b",
    10 => x"80c7c808",
    11 => x"0b0b80c7",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c7cc0c0b",
    16 => x"0b80c7c8",
    17 => x"0c0b0b80",
    18 => x"c7c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb4c0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c7c470",
    57 => x"80d1f427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5189dd",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c7",
    65 => x"d40c9f0b",
    66 => x"80c7d80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c7d808ff",
    70 => x"0580c7d8",
    71 => x"0c80c7d8",
    72 => x"088025e8",
    73 => x"3880c7d4",
    74 => x"08ff0580",
    75 => x"c7d40c80",
    76 => x"c7d40880",
    77 => x"25d03880",
    78 => x"0b80c7d8",
    79 => x"0c800b80",
    80 => x"c7d40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c7d408",
   100 => x"25913882",
   101 => x"c82d80c7",
   102 => x"d408ff05",
   103 => x"80c7d40c",
   104 => x"838a0480",
   105 => x"c7d40880",
   106 => x"c7d80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c7d408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c7d80881",
   116 => x"0580c7d8",
   117 => x"0c80c7d8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c7d8",
   121 => x"0c80c7d4",
   122 => x"08810580",
   123 => x"c7d40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c7",
   128 => x"d8088105",
   129 => x"80c7d80c",
   130 => x"80c7d808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c7d8",
   134 => x"0c80c7d4",
   135 => x"08810580",
   136 => x"c7d40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"c7dc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"c7dc0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280c7",
   177 => x"dc088407",
   178 => x"80c7dc0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b0bbf",
   183 => x"f40c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80c7dc",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80c7",
   208 => x"c40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050d84bf",
   216 => x"5186c72d",
   217 => x"ff115170",
   218 => x"8025f638",
   219 => x"0284050d",
   220 => x"0402fc05",
   221 => x"0dec5183",
   222 => x"710c86c7",
   223 => x"2d82710c",
   224 => x"90c62d02",
   225 => x"84050d04",
   226 => x"02fc050d",
   227 => x"ec518182",
   228 => x"710c86c7",
   229 => x"2d82710c",
   230 => x"90c62d02",
   231 => x"84050d04",
   232 => x"02fc050d",
   233 => x"ec5180c2",
   234 => x"710c86c7",
   235 => x"2d82710c",
   236 => x"90c62d02",
   237 => x"84050d04",
   238 => x"02fc050d",
   239 => x"ec518282",
   240 => x"710c86c7",
   241 => x"2d82710c",
   242 => x"90c62d02",
   243 => x"84050d04",
   244 => x"02fc050d",
   245 => x"ec519271",
   246 => x"0c86c72d",
   247 => x"82710c02",
   248 => x"84050d04",
   249 => x"02d0050d",
   250 => x"7d548074",
   251 => x"5380c7e0",
   252 => x"525babac",
   253 => x"2d80c7c4",
   254 => x"087b2e81",
   255 => x"b63880c7",
   256 => x"e40870f8",
   257 => x"0c891580",
   258 => x"f52d8a16",
   259 => x"80f52d71",
   260 => x"82802905",
   261 => x"881780f5",
   262 => x"2d708480",
   263 => x"802912f4",
   264 => x"0c575556",
   265 => x"58a40bec",
   266 => x"0c7aff19",
   267 => x"585a767b",
   268 => x"2e8b3881",
   269 => x"1a77812a",
   270 => x"585a76f7",
   271 => x"38f71a5a",
   272 => x"815b8078",
   273 => x"2580ec38",
   274 => x"79527651",
   275 => x"84a82d80",
   276 => x"c8ac5280",
   277 => x"c7e051ad",
   278 => x"f92d80c7",
   279 => x"c408802e",
   280 => x"b93880c8",
   281 => x"ac5c83fc",
   282 => x"597b7084",
   283 => x"055d0870",
   284 => x"81ff0671",
   285 => x"882a7081",
   286 => x"ff067390",
   287 => x"2a7081ff",
   288 => x"0675982a",
   289 => x"e80ce80c",
   290 => x"58e80c57",
   291 => x"e80cfc1a",
   292 => x"5a537880",
   293 => x"25d33889",
   294 => x"a20480c7",
   295 => x"c4085b84",
   296 => x"805880c7",
   297 => x"e051adc9",
   298 => x"2dfc8018",
   299 => x"81185858",
   300 => x"88c20486",
   301 => x"da2d840b",
   302 => x"ec0c7a80",
   303 => x"2e8e3880",
   304 => x"c3b45192",
   305 => x"d02d90c6",
   306 => x"2d89d304",
   307 => x"80c59451",
   308 => x"92d02d7a",
   309 => x"80c7c40c",
   310 => x"02b0050d",
   311 => x"0402ec05",
   312 => x"0d840bec",
   313 => x"0c90a42d",
   314 => x"8cf62d81",
   315 => x"f92da1ec",
   316 => x"2d80c7c4",
   317 => x"08802e82",
   318 => x"e63887e4",
   319 => x"51b4b92d",
   320 => x"80c3b451",
   321 => x"92d02d90",
   322 => x"c62d8d82",
   323 => x"2d92e32d",
   324 => x"80c2a80b",
   325 => x"80f52d70",
   326 => x"822b8406",
   327 => x"80c2b40b",
   328 => x"80f52d70",
   329 => x"982b8180",
   330 => x"0a0680c2",
   331 => x"c00b80f5",
   332 => x"2d70842b",
   333 => x"b0067473",
   334 => x"070780c2",
   335 => x"cc0b80f5",
   336 => x"2d70882b",
   337 => x"8e800680",
   338 => x"c2d80b80",
   339 => x"f52d7086",
   340 => x"2b80c006",
   341 => x"74730707",
   342 => x"80c0f00b",
   343 => x"80f52d70",
   344 => x"8d2b80c0",
   345 => x"800680c0",
   346 => x"fc0b80f5",
   347 => x"2d70902b",
   348 => x"84808006",
   349 => x"74730707",
   350 => x"80c1880b",
   351 => x"80f52d70",
   352 => x"942b9c80",
   353 => x"0a0680c1",
   354 => x"940b80f5",
   355 => x"2d708c2b",
   356 => x"a0800674",
   357 => x"73070780",
   358 => x"c1a00b80",
   359 => x"f52d7092",
   360 => x"2bb08080",
   361 => x"0680c1ac",
   362 => x"0b80f52d",
   363 => x"709e2b82",
   364 => x"0a067473",
   365 => x"070780c1",
   366 => x"b80b80f5",
   367 => x"2d709f2b",
   368 => x"720780c0",
   369 => x"800b80f5",
   370 => x"2d70832b",
   371 => x"880680c0",
   372 => x"8c0b80f5",
   373 => x"2d701082",
   374 => x"06747307",
   375 => x"0780c098",
   376 => x"0b80f52d",
   377 => x"709a2bb0",
   378 => x"0a0680c0",
   379 => x"a40b80f5",
   380 => x"2d709c2b",
   381 => x"8c0a0674",
   382 => x"73070780",
   383 => x"c49c0b80",
   384 => x"f52d708e",
   385 => x"2b838080",
   386 => x"0680c4a8",
   387 => x"0b80f52d",
   388 => x"708b2b90",
   389 => x"80067473",
   390 => x"070780c4",
   391 => x"b40b80f5",
   392 => x"2d708106",
   393 => x"a02b7207",
   394 => x"fc0c5354",
   395 => x"54545454",
   396 => x"54545654",
   397 => x"52565452",
   398 => x"54545454",
   399 => x"54545454",
   400 => x"54545454",
   401 => x"54545454",
   402 => x"56545257",
   403 => x"57535386",
   404 => x"5280c7c4",
   405 => x"08833884",
   406 => x"5271ec0c",
   407 => x"8a8a0480",
   408 => x"0b80c7c4",
   409 => x"0c029405",
   410 => x"0d047198",
   411 => x"0c04ffb0",
   412 => x"0880c7c4",
   413 => x"0c04810b",
   414 => x"ffb00c04",
   415 => x"800bffb0",
   416 => x"0c0402f4",
   417 => x"050d8e90",
   418 => x"0480c7c4",
   419 => x"0881f02e",
   420 => x"0981068a",
   421 => x"38810b80",
   422 => x"c5f80c8e",
   423 => x"900480c7",
   424 => x"c40881e0",
   425 => x"2e098106",
   426 => x"8a38810b",
   427 => x"80c5fc0c",
   428 => x"8e900480",
   429 => x"c7c40852",
   430 => x"80c5fc08",
   431 => x"802e8938",
   432 => x"80c7c408",
   433 => x"81800552",
   434 => x"71842c72",
   435 => x"8f065353",
   436 => x"80c5f808",
   437 => x"802e9a38",
   438 => x"72842980",
   439 => x"c5b80572",
   440 => x"1381712b",
   441 => x"70097308",
   442 => x"06730c51",
   443 => x"53538e84",
   444 => x"04728429",
   445 => x"80c5b805",
   446 => x"72138371",
   447 => x"2b720807",
   448 => x"720c5353",
   449 => x"800b80c5",
   450 => x"fc0c800b",
   451 => x"80c5f80c",
   452 => x"80c7ec51",
   453 => x"8f972d80",
   454 => x"c7c408ff",
   455 => x"24feea38",
   456 => x"800b80c7",
   457 => x"c40c028c",
   458 => x"050d0402",
   459 => x"f8050d80",
   460 => x"c5b8528f",
   461 => x"51807270",
   462 => x"8405540c",
   463 => x"ff115170",
   464 => x"8025f238",
   465 => x"0288050d",
   466 => x"0402f005",
   467 => x"0d75518c",
   468 => x"fc2d7082",
   469 => x"2cfc0680",
   470 => x"c5b81172",
   471 => x"109e0671",
   472 => x"0870722a",
   473 => x"70830682",
   474 => x"742b7009",
   475 => x"7406760c",
   476 => x"54515657",
   477 => x"5351538c",
   478 => x"f62d7180",
   479 => x"c7c40c02",
   480 => x"90050d04",
   481 => x"02fc050d",
   482 => x"72518071",
   483 => x"0c800b84",
   484 => x"120c0284",
   485 => x"050d0402",
   486 => x"f0050d75",
   487 => x"70088412",
   488 => x"08535353",
   489 => x"ff547171",
   490 => x"2ea8388c",
   491 => x"fc2d8413",
   492 => x"08708429",
   493 => x"14881170",
   494 => x"087081ff",
   495 => x"06841808",
   496 => x"81118706",
   497 => x"841a0c53",
   498 => x"51555151",
   499 => x"518cf62d",
   500 => x"71547380",
   501 => x"c7c40c02",
   502 => x"90050d04",
   503 => x"02f8050d",
   504 => x"8cfc2de0",
   505 => x"08708b2a",
   506 => x"70810651",
   507 => x"52527080",
   508 => x"2ea13880",
   509 => x"c7ec0870",
   510 => x"842980c7",
   511 => x"f4057381",
   512 => x"ff06710c",
   513 => x"515180c7",
   514 => x"ec088111",
   515 => x"870680c7",
   516 => x"ec0c5180",
   517 => x"0b80c894",
   518 => x"0c8cee2d",
   519 => x"8cf62d02",
   520 => x"88050d04",
   521 => x"02fc050d",
   522 => x"80c7ec51",
   523 => x"8f842d8e",
   524 => x"ab2d8fdc",
   525 => x"518cea2d",
   526 => x"0284050d",
   527 => x"0480c898",
   528 => x"0880c7c4",
   529 => x"0c0402fc",
   530 => x"050d90d0",
   531 => x"048d822d",
   532 => x"80f6518e",
   533 => x"c92d80c7",
   534 => x"c408f238",
   535 => x"80da518e",
   536 => x"c92d80c7",
   537 => x"c408e638",
   538 => x"80c7c408",
   539 => x"80c6840c",
   540 => x"80c7c408",
   541 => x"51858d2d",
   542 => x"0284050d",
   543 => x"0402ec05",
   544 => x"0d765480",
   545 => x"52870b88",
   546 => x"1580f52d",
   547 => x"56537472",
   548 => x"248338a0",
   549 => x"53725183",
   550 => x"842d8112",
   551 => x"8b1580f5",
   552 => x"2d545272",
   553 => x"7225de38",
   554 => x"0294050d",
   555 => x"0402f005",
   556 => x"0d80c898",
   557 => x"085481f9",
   558 => x"2d800b80",
   559 => x"c89c0c73",
   560 => x"08802e81",
   561 => x"8638820b",
   562 => x"80c7d80c",
   563 => x"80c89c08",
   564 => x"8f0680c7",
   565 => x"d40c7308",
   566 => x"5271832e",
   567 => x"96387183",
   568 => x"26893871",
   569 => x"812eaf38",
   570 => x"92b40471",
   571 => x"852e9f38",
   572 => x"92b40488",
   573 => x"1480f52d",
   574 => x"841508be",
   575 => x"c0535452",
   576 => x"86a02d71",
   577 => x"84291370",
   578 => x"08525292",
   579 => x"b8047351",
   580 => x"90fd2d92",
   581 => x"b40480c6",
   582 => x"80088815",
   583 => x"082c7081",
   584 => x"06515271",
   585 => x"802e8738",
   586 => x"bec45192",
   587 => x"b104bec8",
   588 => x"5186a02d",
   589 => x"84140851",
   590 => x"86a02d80",
   591 => x"c89c0881",
   592 => x"0580c89c",
   593 => x"0c8c1454",
   594 => x"91bf0402",
   595 => x"90050d04",
   596 => x"7180c898",
   597 => x"0c91ad2d",
   598 => x"80c89c08",
   599 => x"ff0580c8",
   600 => x"a00c0402",
   601 => x"e8050d80",
   602 => x"c8980880",
   603 => x"c8a40857",
   604 => x"5587518e",
   605 => x"c92d80c7",
   606 => x"c408812a",
   607 => x"70810651",
   608 => x"5271802e",
   609 => x"a338938c",
   610 => x"048d822d",
   611 => x"87518ec9",
   612 => x"2d80c7c4",
   613 => x"08f33880",
   614 => x"c6840881",
   615 => x"327080c6",
   616 => x"840c7052",
   617 => x"52858d2d",
   618 => x"80fe518e",
   619 => x"c92d80c7",
   620 => x"c408802e",
   621 => x"a93880c6",
   622 => x"8408802e",
   623 => x"9238800b",
   624 => x"80c6840c",
   625 => x"8051858d",
   626 => x"2d93cf04",
   627 => x"8d822d80",
   628 => x"fe518ec9",
   629 => x"2d80c7c4",
   630 => x"08f23887",
   631 => x"d02d80c6",
   632 => x"84089038",
   633 => x"81fd518e",
   634 => x"c92d81fa",
   635 => x"518ec92d",
   636 => x"99c80481",
   637 => x"f5518ec9",
   638 => x"2d80c7c4",
   639 => x"08812a70",
   640 => x"81065152",
   641 => x"71802eb3",
   642 => x"3880c8a0",
   643 => x"08527180",
   644 => x"2e8a38ff",
   645 => x"1280c8a0",
   646 => x"0c94bb04",
   647 => x"80c89c08",
   648 => x"1080c89c",
   649 => x"08057084",
   650 => x"29165152",
   651 => x"88120880",
   652 => x"2e8938ff",
   653 => x"51881208",
   654 => x"52712d81",
   655 => x"f2518ec9",
   656 => x"2d80c7c4",
   657 => x"08812a70",
   658 => x"81065152",
   659 => x"71802eb4",
   660 => x"3880c89c",
   661 => x"08ff1180",
   662 => x"c8a00856",
   663 => x"53537372",
   664 => x"258a3881",
   665 => x"1480c8a0",
   666 => x"0c958404",
   667 => x"72101370",
   668 => x"84291651",
   669 => x"52881208",
   670 => x"802e8938",
   671 => x"fe518812",
   672 => x"0852712d",
   673 => x"81fd518e",
   674 => x"c92d80c7",
   675 => x"c408812a",
   676 => x"70810651",
   677 => x"5271802e",
   678 => x"b13880c8",
   679 => x"a008802e",
   680 => x"8a38800b",
   681 => x"80c8a00c",
   682 => x"95ca0480",
   683 => x"c89c0810",
   684 => x"80c89c08",
   685 => x"05708429",
   686 => x"16515288",
   687 => x"1208802e",
   688 => x"8938fd51",
   689 => x"88120852",
   690 => x"712d81fa",
   691 => x"518ec92d",
   692 => x"80c7c408",
   693 => x"812a7081",
   694 => x"06515271",
   695 => x"802eb138",
   696 => x"80c89c08",
   697 => x"ff115452",
   698 => x"80c8a008",
   699 => x"73258938",
   700 => x"7280c8a0",
   701 => x"0c969004",
   702 => x"71101270",
   703 => x"84291651",
   704 => x"52881208",
   705 => x"802e8938",
   706 => x"fc518812",
   707 => x"0852712d",
   708 => x"80c8a008",
   709 => x"70535473",
   710 => x"802e8a38",
   711 => x"8c15ff15",
   712 => x"55559697",
   713 => x"04820b80",
   714 => x"c7d80c71",
   715 => x"8f0680c7",
   716 => x"d40c81eb",
   717 => x"518ec92d",
   718 => x"80c7c408",
   719 => x"812a7081",
   720 => x"06515271",
   721 => x"802ead38",
   722 => x"7408852e",
   723 => x"098106a4",
   724 => x"38881580",
   725 => x"f52dff05",
   726 => x"52718816",
   727 => x"81b72d71",
   728 => x"982b5271",
   729 => x"80258838",
   730 => x"800b8816",
   731 => x"81b72d74",
   732 => x"5190fd2d",
   733 => x"81f4518e",
   734 => x"c92d80c7",
   735 => x"c408812a",
   736 => x"70810651",
   737 => x"5271802e",
   738 => x"b3387408",
   739 => x"852e0981",
   740 => x"06aa3888",
   741 => x"1580f52d",
   742 => x"81055271",
   743 => x"881681b7",
   744 => x"2d7181ff",
   745 => x"068b1680",
   746 => x"f52d5452",
   747 => x"72722787",
   748 => x"38728816",
   749 => x"81b72d74",
   750 => x"5190fd2d",
   751 => x"80da518e",
   752 => x"c92d80c7",
   753 => x"c408812a",
   754 => x"70810651",
   755 => x"5271802e",
   756 => x"81ad3880",
   757 => x"c8980880",
   758 => x"c8a00855",
   759 => x"5373802e",
   760 => x"8a388c13",
   761 => x"ff155553",
   762 => x"97dd0472",
   763 => x"08527182",
   764 => x"2ea63871",
   765 => x"82268938",
   766 => x"71812eaa",
   767 => x"3898ff04",
   768 => x"71832eb4",
   769 => x"3871842e",
   770 => x"09810680",
   771 => x"f2388813",
   772 => x"085192d0",
   773 => x"2d98ff04",
   774 => x"80c8a008",
   775 => x"51881308",
   776 => x"52712d98",
   777 => x"ff04810b",
   778 => x"8814082b",
   779 => x"80c68008",
   780 => x"3280c680",
   781 => x"0c98d304",
   782 => x"881380f5",
   783 => x"2d81058b",
   784 => x"1480f52d",
   785 => x"53547174",
   786 => x"24833880",
   787 => x"54738814",
   788 => x"81b72d91",
   789 => x"ad2d98ff",
   790 => x"04750880",
   791 => x"2ea43875",
   792 => x"08518ec9",
   793 => x"2d80c7c4",
   794 => x"08810652",
   795 => x"71802e8c",
   796 => x"3880c8a0",
   797 => x"08518416",
   798 => x"0852712d",
   799 => x"88165675",
   800 => x"d8388054",
   801 => x"800b80c7",
   802 => x"d80c738f",
   803 => x"0680c7d4",
   804 => x"0ca05273",
   805 => x"80c8a008",
   806 => x"2e098106",
   807 => x"993880c8",
   808 => x"9c08ff05",
   809 => x"74327009",
   810 => x"81057072",
   811 => x"079f2a91",
   812 => x"71315151",
   813 => x"53537151",
   814 => x"83842d81",
   815 => x"14548e74",
   816 => x"25c23880",
   817 => x"c6840852",
   818 => x"7180c7c4",
   819 => x"0c029805",
   820 => x"0d0402f4",
   821 => x"050dd452",
   822 => x"81ff720c",
   823 => x"71085381",
   824 => x"ff720c72",
   825 => x"882b83fe",
   826 => x"80067208",
   827 => x"7081ff06",
   828 => x"51525381",
   829 => x"ff720c72",
   830 => x"7107882b",
   831 => x"72087081",
   832 => x"ff065152",
   833 => x"5381ff72",
   834 => x"0c727107",
   835 => x"882b7208",
   836 => x"7081ff06",
   837 => x"720780c7",
   838 => x"c40c5253",
   839 => x"028c050d",
   840 => x"0402f405",
   841 => x"0d747671",
   842 => x"81ff06d4",
   843 => x"0c535380",
   844 => x"c8a80885",
   845 => x"3871892b",
   846 => x"5271982a",
   847 => x"d40c7190",
   848 => x"2a7081ff",
   849 => x"06d40c51",
   850 => x"71882a70",
   851 => x"81ff06d4",
   852 => x"0c517181",
   853 => x"ff06d40c",
   854 => x"72902a70",
   855 => x"81ff06d4",
   856 => x"0c51d408",
   857 => x"7081ff06",
   858 => x"515182b8",
   859 => x"bf527081",
   860 => x"ff2e0981",
   861 => x"06943881",
   862 => x"ff0bd40c",
   863 => x"d4087081",
   864 => x"ff06ff14",
   865 => x"54515171",
   866 => x"e5387080",
   867 => x"c7c40c02",
   868 => x"8c050d04",
   869 => x"02fc050d",
   870 => x"81c75181",
   871 => x"ff0bd40c",
   872 => x"ff115170",
   873 => x"8025f438",
   874 => x"0284050d",
   875 => x"0402f405",
   876 => x"0d81ff0b",
   877 => x"d40c9353",
   878 => x"805287fc",
   879 => x"80c1519a",
   880 => x"a12d80c7",
   881 => x"c4088b38",
   882 => x"81ff0bd4",
   883 => x"0c81539b",
   884 => x"db049b94",
   885 => x"2dff1353",
   886 => x"72de3872",
   887 => x"80c7c40c",
   888 => x"028c050d",
   889 => x"0402ec05",
   890 => x"0d810b80",
   891 => x"c8a80c84",
   892 => x"54d00870",
   893 => x"8f2a7081",
   894 => x"06515153",
   895 => x"72f33872",
   896 => x"d00c9b94",
   897 => x"2dbecc51",
   898 => x"86a02dd0",
   899 => x"08708f2a",
   900 => x"70810651",
   901 => x"515372f3",
   902 => x"38810bd0",
   903 => x"0cb15380",
   904 => x"5284d480",
   905 => x"c0519aa1",
   906 => x"2d80c7c4",
   907 => x"08812e93",
   908 => x"3872822e",
   909 => x"bf38ff13",
   910 => x"5372e438",
   911 => x"ff145473",
   912 => x"ffaf389b",
   913 => x"942d83aa",
   914 => x"52849c80",
   915 => x"c8519aa1",
   916 => x"2d80c7c4",
   917 => x"08812e09",
   918 => x"81069338",
   919 => x"99d22d80",
   920 => x"c7c40883",
   921 => x"ffff0653",
   922 => x"7283aa2e",
   923 => x"9d389bad",
   924 => x"2d9d8504",
   925 => x"bed85186",
   926 => x"a02d8053",
   927 => x"9eda04be",
   928 => x"f05186a0",
   929 => x"2d80549e",
   930 => x"ab0481ff",
   931 => x"0bd40cb1",
   932 => x"549b942d",
   933 => x"8fcf5380",
   934 => x"5287fc80",
   935 => x"f7519aa1",
   936 => x"2d80c7c4",
   937 => x"085580c7",
   938 => x"c408812e",
   939 => x"0981069c",
   940 => x"3881ff0b",
   941 => x"d40c820a",
   942 => x"52849c80",
   943 => x"e9519aa1",
   944 => x"2d80c7c4",
   945 => x"08802e8d",
   946 => x"389b942d",
   947 => x"ff135372",
   948 => x"c6389e9e",
   949 => x"0481ff0b",
   950 => x"d40c80c7",
   951 => x"c4085287",
   952 => x"fc80fa51",
   953 => x"9aa12d80",
   954 => x"c7c408b2",
   955 => x"3881ff0b",
   956 => x"d40cd408",
   957 => x"5381ff0b",
   958 => x"d40c81ff",
   959 => x"0bd40c81",
   960 => x"ff0bd40c",
   961 => x"81ff0bd4",
   962 => x"0c72862a",
   963 => x"70810676",
   964 => x"56515372",
   965 => x"963880c7",
   966 => x"c408549e",
   967 => x"ab047382",
   968 => x"2efedc38",
   969 => x"ff145473",
   970 => x"fee73873",
   971 => x"80c8a80c",
   972 => x"738b3881",
   973 => x"5287fc80",
   974 => x"d0519aa1",
   975 => x"2d81ff0b",
   976 => x"d40cd008",
   977 => x"708f2a70",
   978 => x"81065151",
   979 => x"5372f338",
   980 => x"72d00c81",
   981 => x"ff0bd40c",
   982 => x"81537280",
   983 => x"c7c40c02",
   984 => x"94050d04",
   985 => x"02e8050d",
   986 => x"78558056",
   987 => x"81ff0bd4",
   988 => x"0cd00870",
   989 => x"8f2a7081",
   990 => x"06515153",
   991 => x"72f33882",
   992 => x"810bd00c",
   993 => x"81ff0bd4",
   994 => x"0c775287",
   995 => x"fc80d151",
   996 => x"9aa12d80",
   997 => x"dbc6df54",
   998 => x"80c7c408",
   999 => x"802e8a38",
  1000 => x"bf905186",
  1001 => x"a02d9ffd",
  1002 => x"0481ff0b",
  1003 => x"d40cd408",
  1004 => x"7081ff06",
  1005 => x"51537281",
  1006 => x"fe2e0981",
  1007 => x"069e3880",
  1008 => x"ff5399d2",
  1009 => x"2d80c7c4",
  1010 => x"08757084",
  1011 => x"05570cff",
  1012 => x"13537280",
  1013 => x"25ec3881",
  1014 => x"569fe204",
  1015 => x"ff145473",
  1016 => x"c83881ff",
  1017 => x"0bd40c81",
  1018 => x"ff0bd40c",
  1019 => x"d008708f",
  1020 => x"2a708106",
  1021 => x"51515372",
  1022 => x"f33872d0",
  1023 => x"0c7580c7",
  1024 => x"c40c0298",
  1025 => x"050d0402",
  1026 => x"e8050d77",
  1027 => x"797b5855",
  1028 => x"55805372",
  1029 => x"7625a338",
  1030 => x"74708105",
  1031 => x"5680f52d",
  1032 => x"74708105",
  1033 => x"5680f52d",
  1034 => x"52527171",
  1035 => x"2e863881",
  1036 => x"51a0bc04",
  1037 => x"811353a0",
  1038 => x"93048051",
  1039 => x"7080c7c4",
  1040 => x"0c029805",
  1041 => x"0d0402ec",
  1042 => x"050d7655",
  1043 => x"74802e80",
  1044 => x"c2389a15",
  1045 => x"80e02d51",
  1046 => x"aed32d80",
  1047 => x"c7c40880",
  1048 => x"c7c40880",
  1049 => x"cedc0c80",
  1050 => x"c7c40854",
  1051 => x"5480ceb8",
  1052 => x"08802e9a",
  1053 => x"38941580",
  1054 => x"e02d51ae",
  1055 => x"d32d80c7",
  1056 => x"c408902b",
  1057 => x"83fff00a",
  1058 => x"06707507",
  1059 => x"51537280",
  1060 => x"cedc0c80",
  1061 => x"cedc0853",
  1062 => x"72802e9d",
  1063 => x"3880ceb0",
  1064 => x"08fe1471",
  1065 => x"2980cec4",
  1066 => x"080580ce",
  1067 => x"e00c7084",
  1068 => x"2b80cebc",
  1069 => x"0c54a1e7",
  1070 => x"0480cec8",
  1071 => x"0880cedc",
  1072 => x"0c80cecc",
  1073 => x"0880cee0",
  1074 => x"0c80ceb8",
  1075 => x"08802e8b",
  1076 => x"3880ceb0",
  1077 => x"08842b53",
  1078 => x"a1e20480",
  1079 => x"ced00884",
  1080 => x"2b537280",
  1081 => x"cebc0c02",
  1082 => x"94050d04",
  1083 => x"02d8050d",
  1084 => x"800b80ce",
  1085 => x"b80c8454",
  1086 => x"9be52d80",
  1087 => x"c7c40880",
  1088 => x"2e973880",
  1089 => x"c8ac5280",
  1090 => x"519ee42d",
  1091 => x"80c7c408",
  1092 => x"802e8638",
  1093 => x"fe54a2a1",
  1094 => x"04ff1454",
  1095 => x"738024d8",
  1096 => x"38738c38",
  1097 => x"bfa05186",
  1098 => x"a02d7355",
  1099 => x"a7ee0480",
  1100 => x"56810b80",
  1101 => x"cee40c88",
  1102 => x"53bfb452",
  1103 => x"80c8e251",
  1104 => x"a0872d80",
  1105 => x"c7c40876",
  1106 => x"2e098106",
  1107 => x"893880c7",
  1108 => x"c40880ce",
  1109 => x"e40c8853",
  1110 => x"bfc05280",
  1111 => x"c8fe51a0",
  1112 => x"872d80c7",
  1113 => x"c4088938",
  1114 => x"80c7c408",
  1115 => x"80cee40c",
  1116 => x"80cee408",
  1117 => x"802e8180",
  1118 => x"3880cbf2",
  1119 => x"0b80f52d",
  1120 => x"80cbf30b",
  1121 => x"80f52d71",
  1122 => x"982b7190",
  1123 => x"2b0780cb",
  1124 => x"f40b80f5",
  1125 => x"2d70882b",
  1126 => x"720780cb",
  1127 => x"f50b80f5",
  1128 => x"2d710780",
  1129 => x"ccaa0b80",
  1130 => x"f52d80cc",
  1131 => x"ab0b80f5",
  1132 => x"2d71882b",
  1133 => x"07535f54",
  1134 => x"525a5657",
  1135 => x"557381ab",
  1136 => x"aa2e0981",
  1137 => x"068e3875",
  1138 => x"51aea22d",
  1139 => x"80c7c408",
  1140 => x"56a3e104",
  1141 => x"7382d4d5",
  1142 => x"2e8738bf",
  1143 => x"cc51a4aa",
  1144 => x"0480c8ac",
  1145 => x"5275519e",
  1146 => x"e42d80c7",
  1147 => x"c4085580",
  1148 => x"c7c40880",
  1149 => x"2e83f738",
  1150 => x"8853bfc0",
  1151 => x"5280c8fe",
  1152 => x"51a0872d",
  1153 => x"80c7c408",
  1154 => x"8a38810b",
  1155 => x"80ceb80c",
  1156 => x"a4b00488",
  1157 => x"53bfb452",
  1158 => x"80c8e251",
  1159 => x"a0872d80",
  1160 => x"c7c40880",
  1161 => x"2e8a38bf",
  1162 => x"e05186a0",
  1163 => x"2da58f04",
  1164 => x"80ccaa0b",
  1165 => x"80f52d54",
  1166 => x"7380d52e",
  1167 => x"09810680",
  1168 => x"ce3880cc",
  1169 => x"ab0b80f5",
  1170 => x"2d547381",
  1171 => x"aa2e0981",
  1172 => x"06bd3880",
  1173 => x"0b80c8ac",
  1174 => x"0b80f52d",
  1175 => x"56547481",
  1176 => x"e92e8338",
  1177 => x"81547481",
  1178 => x"eb2e8c38",
  1179 => x"80557375",
  1180 => x"2e098106",
  1181 => x"82f83880",
  1182 => x"c8b70b80",
  1183 => x"f52d5574",
  1184 => x"8e3880c8",
  1185 => x"b80b80f5",
  1186 => x"2d547382",
  1187 => x"2e863880",
  1188 => x"55a7ee04",
  1189 => x"80c8b90b",
  1190 => x"80f52d70",
  1191 => x"80ceb00c",
  1192 => x"ff0580ce",
  1193 => x"b40c80c8",
  1194 => x"ba0b80f5",
  1195 => x"2d80c8bb",
  1196 => x"0b80f52d",
  1197 => x"58760577",
  1198 => x"82802905",
  1199 => x"7080cec0",
  1200 => x"0c80c8bc",
  1201 => x"0b80f52d",
  1202 => x"7080ced4",
  1203 => x"0c80ceb8",
  1204 => x"08595758",
  1205 => x"76802e81",
  1206 => x"b6388853",
  1207 => x"bfc05280",
  1208 => x"c8fe51a0",
  1209 => x"872d80c7",
  1210 => x"c4088282",
  1211 => x"3880ceb0",
  1212 => x"0870842b",
  1213 => x"80cebc0c",
  1214 => x"7080ced0",
  1215 => x"0c80c8d1",
  1216 => x"0b80f52d",
  1217 => x"80c8d00b",
  1218 => x"80f52d71",
  1219 => x"82802905",
  1220 => x"80c8d20b",
  1221 => x"80f52d70",
  1222 => x"84808029",
  1223 => x"1280c8d3",
  1224 => x"0b80f52d",
  1225 => x"7081800a",
  1226 => x"29127080",
  1227 => x"ced80c80",
  1228 => x"ced40871",
  1229 => x"2980cec0",
  1230 => x"08057080",
  1231 => x"cec40c80",
  1232 => x"c8d90b80",
  1233 => x"f52d80c8",
  1234 => x"d80b80f5",
  1235 => x"2d718280",
  1236 => x"290580c8",
  1237 => x"da0b80f5",
  1238 => x"2d708480",
  1239 => x"80291280",
  1240 => x"c8db0b80",
  1241 => x"f52d7098",
  1242 => x"2b81f00a",
  1243 => x"06720570",
  1244 => x"80cec80c",
  1245 => x"fe117e29",
  1246 => x"770580ce",
  1247 => x"cc0c5259",
  1248 => x"5243545e",
  1249 => x"51525952",
  1250 => x"5d575957",
  1251 => x"a7e70480",
  1252 => x"c8be0b80",
  1253 => x"f52d80c8",
  1254 => x"bd0b80f5",
  1255 => x"2d718280",
  1256 => x"29057080",
  1257 => x"cebc0c70",
  1258 => x"a02983ff",
  1259 => x"0570892a",
  1260 => x"7080ced0",
  1261 => x"0c80c8c3",
  1262 => x"0b80f52d",
  1263 => x"80c8c20b",
  1264 => x"80f52d71",
  1265 => x"82802905",
  1266 => x"7080ced8",
  1267 => x"0c7b7129",
  1268 => x"1e7080ce",
  1269 => x"cc0c7d80",
  1270 => x"cec80c73",
  1271 => x"0580cec4",
  1272 => x"0c555e51",
  1273 => x"51555580",
  1274 => x"51a0c62d",
  1275 => x"81557480",
  1276 => x"c7c40c02",
  1277 => x"a8050d04",
  1278 => x"02ec050d",
  1279 => x"7670872c",
  1280 => x"7180ff06",
  1281 => x"55565480",
  1282 => x"ceb8088a",
  1283 => x"3873882c",
  1284 => x"7481ff06",
  1285 => x"545580c8",
  1286 => x"ac5280ce",
  1287 => x"c0081551",
  1288 => x"9ee42d80",
  1289 => x"c7c40854",
  1290 => x"80c7c408",
  1291 => x"802eb838",
  1292 => x"80ceb808",
  1293 => x"802e9a38",
  1294 => x"72842980",
  1295 => x"c8ac0570",
  1296 => x"085253ae",
  1297 => x"a22d80c7",
  1298 => x"c408f00a",
  1299 => x"0653a8e5",
  1300 => x"04721080",
  1301 => x"c8ac0570",
  1302 => x"80e02d52",
  1303 => x"53aed32d",
  1304 => x"80c7c408",
  1305 => x"53725473",
  1306 => x"80c7c40c",
  1307 => x"0294050d",
  1308 => x"0402e005",
  1309 => x"0d797084",
  1310 => x"2c80cee0",
  1311 => x"0805718f",
  1312 => x"06525553",
  1313 => x"728a3880",
  1314 => x"c8ac5273",
  1315 => x"519ee42d",
  1316 => x"72a02980",
  1317 => x"c8ac0554",
  1318 => x"807480f5",
  1319 => x"2d565374",
  1320 => x"732e8338",
  1321 => x"81537481",
  1322 => x"e52e81f4",
  1323 => x"38817074",
  1324 => x"06545872",
  1325 => x"802e81e8",
  1326 => x"388b1480",
  1327 => x"f52d7083",
  1328 => x"2a790658",
  1329 => x"56769b38",
  1330 => x"80c68808",
  1331 => x"53728938",
  1332 => x"7280ccac",
  1333 => x"0b81b72d",
  1334 => x"7680c688",
  1335 => x"0c7353ab",
  1336 => x"a204758f",
  1337 => x"2e098106",
  1338 => x"81b63874",
  1339 => x"9f068d29",
  1340 => x"80cc9f11",
  1341 => x"51538114",
  1342 => x"80f52d73",
  1343 => x"70810555",
  1344 => x"81b72d83",
  1345 => x"1480f52d",
  1346 => x"73708105",
  1347 => x"5581b72d",
  1348 => x"851480f5",
  1349 => x"2d737081",
  1350 => x"055581b7",
  1351 => x"2d871480",
  1352 => x"f52d7370",
  1353 => x"81055581",
  1354 => x"b72d8914",
  1355 => x"80f52d73",
  1356 => x"70810555",
  1357 => x"81b72d8e",
  1358 => x"1480f52d",
  1359 => x"73708105",
  1360 => x"5581b72d",
  1361 => x"901480f5",
  1362 => x"2d737081",
  1363 => x"055581b7",
  1364 => x"2d921480",
  1365 => x"f52d7370",
  1366 => x"81055581",
  1367 => x"b72d9414",
  1368 => x"80f52d73",
  1369 => x"70810555",
  1370 => x"81b72d96",
  1371 => x"1480f52d",
  1372 => x"73708105",
  1373 => x"5581b72d",
  1374 => x"981480f5",
  1375 => x"2d737081",
  1376 => x"055581b7",
  1377 => x"2d9c1480",
  1378 => x"f52d7370",
  1379 => x"81055581",
  1380 => x"b72d9e14",
  1381 => x"80f52d73",
  1382 => x"81b72d77",
  1383 => x"80c6880c",
  1384 => x"80537280",
  1385 => x"c7c40c02",
  1386 => x"a0050d04",
  1387 => x"02cc050d",
  1388 => x"7e605e5a",
  1389 => x"800b80ce",
  1390 => x"dc0880ce",
  1391 => x"e008595c",
  1392 => x"56805880",
  1393 => x"cebc0878",
  1394 => x"2e81b838",
  1395 => x"778f06a0",
  1396 => x"17575473",
  1397 => x"913880c8",
  1398 => x"ac527651",
  1399 => x"8117579e",
  1400 => x"e42d80c8",
  1401 => x"ac568076",
  1402 => x"80f52d56",
  1403 => x"5474742e",
  1404 => x"83388154",
  1405 => x"7481e52e",
  1406 => x"80fd3881",
  1407 => x"70750655",
  1408 => x"5c73802e",
  1409 => x"80f1388b",
  1410 => x"1680f52d",
  1411 => x"98065978",
  1412 => x"80e5388b",
  1413 => x"537c5275",
  1414 => x"51a0872d",
  1415 => x"80c7c408",
  1416 => x"80d5389c",
  1417 => x"160851ae",
  1418 => x"a22d80c7",
  1419 => x"c408841b",
  1420 => x"0c9a1680",
  1421 => x"e02d51ae",
  1422 => x"d32d80c7",
  1423 => x"c40880c7",
  1424 => x"c408881c",
  1425 => x"0c80c7c4",
  1426 => x"08555580",
  1427 => x"ceb80880",
  1428 => x"2e993894",
  1429 => x"1680e02d",
  1430 => x"51aed32d",
  1431 => x"80c7c408",
  1432 => x"902b83ff",
  1433 => x"f00a0670",
  1434 => x"16515473",
  1435 => x"881b0c78",
  1436 => x"7a0c7b54",
  1437 => x"adbf0481",
  1438 => x"185880ce",
  1439 => x"bc087826",
  1440 => x"feca3880",
  1441 => x"ceb80880",
  1442 => x"2eb3387a",
  1443 => x"51a7f82d",
  1444 => x"80c7c408",
  1445 => x"80c7c408",
  1446 => x"80ffffff",
  1447 => x"f806555b",
  1448 => x"7380ffff",
  1449 => x"fff82e95",
  1450 => x"3880c7c4",
  1451 => x"08fe0580",
  1452 => x"ceb00829",
  1453 => x"80cec408",
  1454 => x"0557abc1",
  1455 => x"04805473",
  1456 => x"80c7c40c",
  1457 => x"02b4050d",
  1458 => x"0402f405",
  1459 => x"0d747008",
  1460 => x"8105710c",
  1461 => x"700880ce",
  1462 => x"b4080653",
  1463 => x"53718f38",
  1464 => x"88130851",
  1465 => x"a7f82d80",
  1466 => x"c7c40888",
  1467 => x"140c810b",
  1468 => x"80c7c40c",
  1469 => x"028c050d",
  1470 => x"0402f005",
  1471 => x"0d758811",
  1472 => x"08fe0580",
  1473 => x"ceb00829",
  1474 => x"80cec408",
  1475 => x"11720880",
  1476 => x"ceb40806",
  1477 => x"05795553",
  1478 => x"54549ee4",
  1479 => x"2d029005",
  1480 => x"0d0402f4",
  1481 => x"050d7470",
  1482 => x"882a83fe",
  1483 => x"80067072",
  1484 => x"982a0772",
  1485 => x"882b87fc",
  1486 => x"80800673",
  1487 => x"982b81f0",
  1488 => x"0a067173",
  1489 => x"070780c7",
  1490 => x"c40c5651",
  1491 => x"5351028c",
  1492 => x"050d0402",
  1493 => x"f8050d02",
  1494 => x"8e0580f5",
  1495 => x"2d74882b",
  1496 => x"077083ff",
  1497 => x"ff0680c7",
  1498 => x"c40c5102",
  1499 => x"88050d04",
  1500 => x"02f4050d",
  1501 => x"74767853",
  1502 => x"54528071",
  1503 => x"25973872",
  1504 => x"70810554",
  1505 => x"80f52d72",
  1506 => x"70810554",
  1507 => x"81b72dff",
  1508 => x"115170eb",
  1509 => x"38807281",
  1510 => x"b72d028c",
  1511 => x"050d0402",
  1512 => x"e8050d77",
  1513 => x"56807056",
  1514 => x"54737624",
  1515 => x"b63880ce",
  1516 => x"bc08742e",
  1517 => x"ae387351",
  1518 => x"a8f12d80",
  1519 => x"c7c40880",
  1520 => x"c7c40809",
  1521 => x"81057080",
  1522 => x"c7c40807",
  1523 => x"9f2a7705",
  1524 => x"81175757",
  1525 => x"53537476",
  1526 => x"24893880",
  1527 => x"cebc0874",
  1528 => x"26d43872",
  1529 => x"80c7c40c",
  1530 => x"0298050d",
  1531 => x"0402f005",
  1532 => x"0d80c7c0",
  1533 => x"081651af",
  1534 => x"9f2d80c7",
  1535 => x"c408802e",
  1536 => x"9f388b53",
  1537 => x"80c7c408",
  1538 => x"5280ccac",
  1539 => x"51aef02d",
  1540 => x"80cee808",
  1541 => x"5473802e",
  1542 => x"873880cc",
  1543 => x"ac51732d",
  1544 => x"0290050d",
  1545 => x"0402dc05",
  1546 => x"0d80705a",
  1547 => x"557480c7",
  1548 => x"c00825b4",
  1549 => x"3880cebc",
  1550 => x"08752eac",
  1551 => x"387851a8",
  1552 => x"f12d80c7",
  1553 => x"c4080981",
  1554 => x"057080c7",
  1555 => x"c408079f",
  1556 => x"2a760581",
  1557 => x"1b5b5654",
  1558 => x"7480c7c0",
  1559 => x"08258938",
  1560 => x"80cebc08",
  1561 => x"7926d638",
  1562 => x"80557880",
  1563 => x"cebc0827",
  1564 => x"81db3878",
  1565 => x"51a8f12d",
  1566 => x"80c7c408",
  1567 => x"802e81ad",
  1568 => x"3880c7c4",
  1569 => x"088b0580",
  1570 => x"f52d7084",
  1571 => x"2a708106",
  1572 => x"77107884",
  1573 => x"2b80ccac",
  1574 => x"0b80f52d",
  1575 => x"5c5c5351",
  1576 => x"55567380",
  1577 => x"2e80cb38",
  1578 => x"7416822b",
  1579 => x"b2f10b80",
  1580 => x"c694120c",
  1581 => x"54777531",
  1582 => x"1080ceec",
  1583 => x"11555690",
  1584 => x"74708105",
  1585 => x"5681b72d",
  1586 => x"a07481b7",
  1587 => x"2d7681ff",
  1588 => x"06811658",
  1589 => x"5473802e",
  1590 => x"8a389c53",
  1591 => x"80ccac52",
  1592 => x"b1ea048b",
  1593 => x"5380c7c4",
  1594 => x"085280ce",
  1595 => x"ee1651b2",
  1596 => x"a5047416",
  1597 => x"822bafed",
  1598 => x"0b80c694",
  1599 => x"120c5476",
  1600 => x"81ff0681",
  1601 => x"16585473",
  1602 => x"802e8a38",
  1603 => x"9c5380cc",
  1604 => x"ac52b29c",
  1605 => x"048b5380",
  1606 => x"c7c40852",
  1607 => x"77753110",
  1608 => x"80ceec05",
  1609 => x"517655ae",
  1610 => x"f02db2c2",
  1611 => x"04749029",
  1612 => x"75317010",
  1613 => x"80ceec05",
  1614 => x"515480c7",
  1615 => x"c4087481",
  1616 => x"b72d8119",
  1617 => x"59748b24",
  1618 => x"a338b0ea",
  1619 => x"04749029",
  1620 => x"75317010",
  1621 => x"80ceec05",
  1622 => x"8c773157",
  1623 => x"51548074",
  1624 => x"81b72d9e",
  1625 => x"14ff1656",
  1626 => x"5474f338",
  1627 => x"02a4050d",
  1628 => x"0402fc05",
  1629 => x"0d80c7c0",
  1630 => x"081351af",
  1631 => x"9f2d80c7",
  1632 => x"c408802e",
  1633 => x"893880c7",
  1634 => x"c40851a0",
  1635 => x"c62d800b",
  1636 => x"80c7c00c",
  1637 => x"b0a52d91",
  1638 => x"ad2d0284",
  1639 => x"050d0402",
  1640 => x"fc050d72",
  1641 => x"5170fd2e",
  1642 => x"b03870fd",
  1643 => x"248a3870",
  1644 => x"fc2e80cc",
  1645 => x"38b48a04",
  1646 => x"70fe2eb7",
  1647 => x"3870ff2e",
  1648 => x"09810680",
  1649 => x"c53880c7",
  1650 => x"c0085170",
  1651 => x"802ebb38",
  1652 => x"ff1180c7",
  1653 => x"c00cb48a",
  1654 => x"0480c7c0",
  1655 => x"08f00570",
  1656 => x"80c7c00c",
  1657 => x"51708025",
  1658 => x"a138800b",
  1659 => x"80c7c00c",
  1660 => x"b48a0480",
  1661 => x"c7c00881",
  1662 => x"0580c7c0",
  1663 => x"0cb48a04",
  1664 => x"80c7c008",
  1665 => x"900580c7",
  1666 => x"c00cb0a5",
  1667 => x"2d91ad2d",
  1668 => x"0284050d",
  1669 => x"0402fc05",
  1670 => x"0d800b80",
  1671 => x"c7c00cb0",
  1672 => x"a52d90bd",
  1673 => x"2d80c7c4",
  1674 => x"0880c7b0",
  1675 => x"0c80c68c",
  1676 => x"5192d02d",
  1677 => x"0284050d",
  1678 => x"047180ce",
  1679 => x"e80c0400",
  1680 => x"00ffffff",
  1681 => x"ff00ffff",
  1682 => x"ffff00ff",
  1683 => x"ffffff00",
  1684 => x"45786974",
  1685 => x"00000000",
  1686 => x"506f7420",
  1687 => x"33263420",
  1688 => x"4a6f7920",
  1689 => x"32204469",
  1690 => x"73706172",
  1691 => x"6f20322f",
  1692 => x"33000000",
  1693 => x"506f7420",
  1694 => x"33263420",
  1695 => x"5261746f",
  1696 => x"6e000000",
  1697 => x"506f7420",
  1698 => x"33263420",
  1699 => x"50616464",
  1700 => x"6c657320",
  1701 => x"33263400",
  1702 => x"506f7420",
  1703 => x"31263220",
  1704 => x"4a6f7920",
  1705 => x"31204469",
  1706 => x"73706172",
  1707 => x"6f20322f",
  1708 => x"33000000",
  1709 => x"506f7420",
  1710 => x"31263220",
  1711 => x"5261746f",
  1712 => x"6e000000",
  1713 => x"506f7420",
  1714 => x"31263220",
  1715 => x"50616464",
  1716 => x"6c657320",
  1717 => x"31263200",
  1718 => x"50756572",
  1719 => x"746f2055",
  1720 => x"41525400",
  1721 => x"50756572",
  1722 => x"746f204a",
  1723 => x"6f797374",
  1724 => x"69636b73",
  1725 => x"00000000",
  1726 => x"4a6f7973",
  1727 => x"7469636b",
  1728 => x"73204e6f",
  1729 => x"726d616c",
  1730 => x"00000000",
  1731 => x"4a6f7973",
  1732 => x"7469636b",
  1733 => x"7320496e",
  1734 => x"74657263",
  1735 => x"616d6269",
  1736 => x"61646f73",
  1737 => x"00000000",
  1738 => x"53696420",
  1739 => x"64696769",
  1740 => x"74616c20",
  1741 => x"61204469",
  1742 => x"67696d61",
  1743 => x"78204e6f",
  1744 => x"00000000",
  1745 => x"53696420",
  1746 => x"64696769",
  1747 => x"74616c20",
  1748 => x"61204469",
  1749 => x"67696d61",
  1750 => x"78205369",
  1751 => x"00000000",
  1752 => x"44696769",
  1753 => x"6d617820",
  1754 => x"4e6f0000",
  1755 => x"44696769",
  1756 => x"6d617820",
  1757 => x"53690000",
  1758 => x"4d657a63",
  1759 => x"6c612053",
  1760 => x"74657265",
  1761 => x"6f204e6f",
  1762 => x"00000000",
  1763 => x"4d657a63",
  1764 => x"6c612053",
  1765 => x"74657265",
  1766 => x"6f203235",
  1767 => x"25000000",
  1768 => x"4d657a63",
  1769 => x"6c612053",
  1770 => x"74657265",
  1771 => x"6f203530",
  1772 => x"25000000",
  1773 => x"4d657a63",
  1774 => x"6c612053",
  1775 => x"74657265",
  1776 => x"6f203735",
  1777 => x"25000000",
  1778 => x"45787061",
  1779 => x"6e73696f",
  1780 => x"6e206465",
  1781 => x"20536f6e",
  1782 => x"69646f20",
  1783 => x"4e6f0000",
  1784 => x"45787061",
  1785 => x"6e73696f",
  1786 => x"6e206465",
  1787 => x"20536f6e",
  1788 => x"69646f20",
  1789 => x"4f504c32",
  1790 => x"00000000",
  1791 => x"53494420",
  1792 => x"44657265",
  1793 => x"63686f20",
  1794 => x"41646472",
  1795 => x"20496775",
  1796 => x"616c0000",
  1797 => x"53494420",
  1798 => x"44657265",
  1799 => x"63686f20",
  1800 => x"41646472",
  1801 => x"20444530",
  1802 => x"30000000",
  1803 => x"53494420",
  1804 => x"44657265",
  1805 => x"63686f20",
  1806 => x"41646472",
  1807 => x"20443432",
  1808 => x"30000000",
  1809 => x"53494420",
  1810 => x"44657265",
  1811 => x"63686f20",
  1812 => x"41646472",
  1813 => x"20443530",
  1814 => x"30000000",
  1815 => x"53494420",
  1816 => x"44657265",
  1817 => x"63686f20",
  1818 => x"41646472",
  1819 => x"20444630",
  1820 => x"30000000",
  1821 => x"53494420",
  1822 => x"44657265",
  1823 => x"63686f20",
  1824 => x"36353831",
  1825 => x"00000000",
  1826 => x"53494420",
  1827 => x"44657265",
  1828 => x"63686f20",
  1829 => x"38353830",
  1830 => x"00000000",
  1831 => x"53494420",
  1832 => x"497a7175",
  1833 => x"69657264",
  1834 => x"6f203635",
  1835 => x"38310000",
  1836 => x"53494420",
  1837 => x"497a7175",
  1838 => x"69657264",
  1839 => x"6f203835",
  1840 => x"38300000",
  1841 => x"50616c65",
  1842 => x"74612043",
  1843 => x"36340000",
  1844 => x"50616c65",
  1845 => x"74612043",
  1846 => x"65506543",
  1847 => x"65526100",
  1848 => x"5363616e",
  1849 => x"646f7562",
  1850 => x"6c657220",
  1851 => x"4e696e67",
  1852 => x"756e6f00",
  1853 => x"5363616e",
  1854 => x"646f7562",
  1855 => x"6c657220",
  1856 => x"48513278",
  1857 => x"2d333230",
  1858 => x"00000000",
  1859 => x"5363616e",
  1860 => x"646f7562",
  1861 => x"6c657220",
  1862 => x"48513278",
  1863 => x"2d313630",
  1864 => x"00000000",
  1865 => x"5363616e",
  1866 => x"646f7562",
  1867 => x"6c657220",
  1868 => x"43525420",
  1869 => x"32352500",
  1870 => x"5363616e",
  1871 => x"646f7562",
  1872 => x"6c657220",
  1873 => x"43525420",
  1874 => x"35302500",
  1875 => x"5363616e",
  1876 => x"646f7562",
  1877 => x"6c657220",
  1878 => x"43525420",
  1879 => x"37352500",
  1880 => x"466f726d",
  1881 => x"61746f20",
  1882 => x"4f726967",
  1883 => x"696e616c",
  1884 => x"00000000",
  1885 => x"466f726d",
  1886 => x"61746f20",
  1887 => x"50616e74",
  1888 => x"616c6c61",
  1889 => x"20436f6d",
  1890 => x"706c6574",
  1891 => x"61000000",
  1892 => x"466f726d",
  1893 => x"61746f20",
  1894 => x"5b415243",
  1895 => x"315d0000",
  1896 => x"466f726d",
  1897 => x"61746f20",
  1898 => x"5b415243",
  1899 => x"325d0000",
  1900 => x"41737065",
  1901 => x"63746f20",
  1902 => x"4f726967",
  1903 => x"696e616c",
  1904 => x"00000000",
  1905 => x"41737065",
  1906 => x"63746f20",
  1907 => x"416e6368",
  1908 => x"6f000000",
  1909 => x"56696465",
  1910 => x"6f205041",
  1911 => x"4c000000",
  1912 => x"56696465",
  1913 => x"6f204e54",
  1914 => x"53430000",
  1915 => x"2020203d",
  1916 => x"20434f4d",
  1917 => x"4f444f52",
  1918 => x"45202036",
  1919 => x"34203d20",
  1920 => x"20200000",
  1921 => x"20202020",
  1922 => x"20204e65",
  1923 => x"75726f52",
  1924 => x"756c657a",
  1925 => x"20202020",
  1926 => x"20200000",
  1927 => x"20202020",
  1928 => x"20202020",
  1929 => x"20202020",
  1930 => x"20202020",
  1931 => x"20202020",
  1932 => x"20200000",
  1933 => x"52657365",
  1934 => x"74000000",
  1935 => x"52657365",
  1936 => x"74202620",
  1937 => x"536f6c74",
  1938 => x"61722043",
  1939 => x"61727475",
  1940 => x"63686f00",
  1941 => x"56696465",
  1942 => x"6f201000",
  1943 => x"41756469",
  1944 => x"6f201000",
  1945 => x"50756572",
  1946 => x"746f7320",
  1947 => x"10000000",
  1948 => x"53616361",
  1949 => x"72204369",
  1950 => x"6e746100",
  1951 => x"506c6179",
  1952 => x"2f53746f",
  1953 => x"70204369",
  1954 => x"6e746100",
  1955 => x"43617267",
  1956 => x"61722044",
  1957 => x"6973636f",
  1958 => x"2f43696e",
  1959 => x"74612f43",
  1960 => x"61727420",
  1961 => x"10000000",
  1962 => x"44697363",
  1963 => x"6f204772",
  1964 => x"61626162",
  1965 => x"6c650000",
  1966 => x"44697363",
  1967 => x"6f20536f",
  1968 => x"6c6f204c",
  1969 => x"65637475",
  1970 => x"72610000",
  1971 => x"536f6e69",
  1972 => x"646f2043",
  1973 => x"696e7461",
  1974 => x"204f6666",
  1975 => x"00000000",
  1976 => x"536f6e69",
  1977 => x"646f2043",
  1978 => x"696e7461",
  1979 => x"204f6e00",
  1980 => x"4b65726e",
  1981 => x"656c2043",
  1982 => x"61726761",
  1983 => x"626c6500",
  1984 => x"4b65726e",
  1985 => x"656c2043",
  1986 => x"36340000",
  1987 => x"4b65726e",
  1988 => x"656c2043",
  1989 => x"36344753",
  1990 => x"00000000",
  1991 => x"4b65726e",
  1992 => x"656c204a",
  1993 => x"61706f6e",
  1994 => x"65730000",
  1995 => x"43617267",
  1996 => x"61204661",
  1997 => x"6c6c6964",
  1998 => x"61000000",
  1999 => x"4f4b0000",
  2000 => x"16200000",
  2001 => x"14200000",
  2002 => x"15200000",
  2003 => x"53442069",
  2004 => x"6e69742e",
  2005 => x"2e2e0a00",
  2006 => x"53442063",
  2007 => x"61726420",
  2008 => x"72657365",
  2009 => x"74206661",
  2010 => x"696c6564",
  2011 => x"210a0000",
  2012 => x"53444843",
  2013 => x"20657272",
  2014 => x"6f72210a",
  2015 => x"00000000",
  2016 => x"57726974",
  2017 => x"65206661",
  2018 => x"696c6564",
  2019 => x"0a000000",
  2020 => x"52656164",
  2021 => x"20666169",
  2022 => x"6c65640a",
  2023 => x"00000000",
  2024 => x"43617264",
  2025 => x"20696e69",
  2026 => x"74206661",
  2027 => x"696c6564",
  2028 => x"0a000000",
  2029 => x"46415431",
  2030 => x"36202020",
  2031 => x"00000000",
  2032 => x"46415433",
  2033 => x"32202020",
  2034 => x"00000000",
  2035 => x"4e6f2070",
  2036 => x"61727469",
  2037 => x"74696f6e",
  2038 => x"20736967",
  2039 => x"0a000000",
  2040 => x"42616420",
  2041 => x"70617274",
  2042 => x"0a000000",
  2043 => x"4261636b",
  2044 => x"00000000",
  2045 => x"00000002",
  2046 => x"00000003",
  2047 => x"00002060",
  2048 => x"00000002",
  2049 => x"00000003",
  2050 => x"00002058",
  2051 => x"00000002",
  2052 => x"00000003",
  2053 => x"0000204c",
  2054 => x"00000003",
  2055 => x"00000003",
  2056 => x"00002040",
  2057 => x"00000003",
  2058 => x"00000004",
  2059 => x"00001a50",
  2060 => x"000021b4",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00001a58",
  2065 => x"00001a74",
  2066 => x"00001a84",
  2067 => x"00001a98",
  2068 => x"00001ab4",
  2069 => x"00001ac4",
  2070 => x"00001ad8",
  2071 => x"00001ae4",
  2072 => x"00001af8",
  2073 => x"00001b0c",
  2074 => x"00000003",
  2075 => x"00002118",
  2076 => x"00000002",
  2077 => x"00000003",
  2078 => x"00002110",
  2079 => x"00000002",
  2080 => x"00000003",
  2081 => x"000020fc",
  2082 => x"00000005",
  2083 => x"00000003",
  2084 => x"000020f4",
  2085 => x"00000002",
  2086 => x"00000003",
  2087 => x"000020e4",
  2088 => x"00000004",
  2089 => x"00000003",
  2090 => x"000020dc",
  2091 => x"00000002",
  2092 => x"00000003",
  2093 => x"000020d4",
  2094 => x"00000002",
  2095 => x"00000004",
  2096 => x"00001a50",
  2097 => x"000021b4",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00001b28",
  2102 => x"00001b44",
  2103 => x"00001b60",
  2104 => x"00001b6c",
  2105 => x"00001b78",
  2106 => x"00001b8c",
  2107 => x"00001ba0",
  2108 => x"00001bb4",
  2109 => x"00001bc8",
  2110 => x"00001be0",
  2111 => x"00001bfc",
  2112 => x"00001c14",
  2113 => x"00001c2c",
  2114 => x"00001c44",
  2115 => x"00001c5c",
  2116 => x"00001c74",
  2117 => x"00001c88",
  2118 => x"00001c9c",
  2119 => x"00001cb0",
  2120 => x"00000003",
  2121 => x"000021ac",
  2122 => x"00000002",
  2123 => x"00000003",
  2124 => x"000021a4",
  2125 => x"00000002",
  2126 => x"00000003",
  2127 => x"00002194",
  2128 => x"00000004",
  2129 => x"00000003",
  2130 => x"0000217c",
  2131 => x"00000006",
  2132 => x"00000003",
  2133 => x"00002174",
  2134 => x"00000002",
  2135 => x"00000004",
  2136 => x"00001a50",
  2137 => x"000021b4",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00001cc4",
  2142 => x"00001cd0",
  2143 => x"00001ce0",
  2144 => x"00001cf4",
  2145 => x"00001d0c",
  2146 => x"00001d24",
  2147 => x"00001d38",
  2148 => x"00001d4c",
  2149 => x"00001d60",
  2150 => x"00001d74",
  2151 => x"00001d90",
  2152 => x"00001da0",
  2153 => x"00001db0",
  2154 => x"00001dc4",
  2155 => x"00001dd4",
  2156 => x"00001de0",
  2157 => x"00000002",
  2158 => x"00001dec",
  2159 => x"00000000",
  2160 => x"00000002",
  2161 => x"00001e04",
  2162 => x"00000000",
  2163 => x"00000002",
  2164 => x"00001e1c",
  2165 => x"00000000",
  2166 => x"00000002",
  2167 => x"00001e34",
  2168 => x"00000371",
  2169 => x"00000002",
  2170 => x"00001e3c",
  2171 => x"00000388",
  2172 => x"00000004",
  2173 => x"00001e54",
  2174 => x"00002120",
  2175 => x"00000004",
  2176 => x"00001e5c",
  2177 => x"00002068",
  2178 => x"00000004",
  2179 => x"00001e64",
  2180 => x"00001ff8",
  2181 => x"00000003",
  2182 => x"00002284",
  2183 => x"00000004",
  2184 => x"00000003",
  2185 => x"0000227c",
  2186 => x"00000002",
  2187 => x"00000003",
  2188 => x"00002274",
  2189 => x"00000002",
  2190 => x"00000002",
  2191 => x"00001e70",
  2192 => x"000003b8",
  2193 => x"00000002",
  2194 => x"00001e7c",
  2195 => x"000003a0",
  2196 => x"00000002",
  2197 => x"00001e8c",
  2198 => x"00001a15",
  2199 => x"00000002",
  2200 => x"00001a50",
  2201 => x"00000846",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00001ea8",
  2206 => x"00001eb8",
  2207 => x"00001ecc",
  2208 => x"00001ee0",
  2209 => x"00001ef0",
  2210 => x"00001f00",
  2211 => x"00001f0c",
  2212 => x"00001f1c",
  2213 => x"00000004",
  2214 => x"00001f2c",
  2215 => x"00002294",
  2216 => x"00000004",
  2217 => x"00001f3c",
  2218 => x"000021b4",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000002",
  2244 => x"0000276c",
  2245 => x"000017ed",
  2246 => x"00000002",
  2247 => x"0000278a",
  2248 => x"000017ed",
  2249 => x"00000002",
  2250 => x"000027a8",
  2251 => x"000017ed",
  2252 => x"00000002",
  2253 => x"000027c6",
  2254 => x"000017ed",
  2255 => x"00000002",
  2256 => x"000027e4",
  2257 => x"000017ed",
  2258 => x"00000002",
  2259 => x"00002802",
  2260 => x"000017ed",
  2261 => x"00000002",
  2262 => x"00002820",
  2263 => x"000017ed",
  2264 => x"00000002",
  2265 => x"0000283e",
  2266 => x"000017ed",
  2267 => x"00000002",
  2268 => x"0000285c",
  2269 => x"000017ed",
  2270 => x"00000002",
  2271 => x"0000287a",
  2272 => x"000017ed",
  2273 => x"00000002",
  2274 => x"00002898",
  2275 => x"000017ed",
  2276 => x"00000002",
  2277 => x"000028b6",
  2278 => x"000017ed",
  2279 => x"00000002",
  2280 => x"000028d4",
  2281 => x"000017ed",
  2282 => x"00000004",
  2283 => x"00001fec",
  2284 => x"00000000",
  2285 => x"00000000",
  2286 => x"00000000",
  2287 => x"0000199f",
  2288 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

