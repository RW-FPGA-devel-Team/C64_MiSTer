-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c6",
     9 => x"b8080b0b",
    10 => x"80c6bc08",
    11 => x"0b0b80c6",
    12 => x"c0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c6c00c0b",
    16 => x"0b80c6bc",
    17 => x"0c0b0b80",
    18 => x"c6b80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb4a0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c6b870",
    57 => x"80d0e827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5189dd",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c6",
    65 => x"c80c9f0b",
    66 => x"80c6cc0c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c6cc08ff",
    70 => x"0580c6cc",
    71 => x"0c80c6cc",
    72 => x"088025e8",
    73 => x"3880c6c8",
    74 => x"08ff0580",
    75 => x"c6c80c80",
    76 => x"c6c80880",
    77 => x"25d03880",
    78 => x"0b80c6cc",
    79 => x"0c800b80",
    80 => x"c6c80c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c6c808",
   100 => x"25913882",
   101 => x"c82d80c6",
   102 => x"c808ff05",
   103 => x"80c6c80c",
   104 => x"838a0480",
   105 => x"c6c80880",
   106 => x"c6cc0853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c6c808",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c6cc0881",
   116 => x"0580c6cc",
   117 => x"0c80c6cc",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c6cc",
   121 => x"0c80c6c8",
   122 => x"08810580",
   123 => x"c6c80c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c6",
   128 => x"cc088105",
   129 => x"80c6cc0c",
   130 => x"80c6cc08",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c6cc",
   134 => x"0c80c6c8",
   135 => x"08810580",
   136 => x"c6c80c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"c6d00cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"c6d00c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280c6",
   177 => x"d0088407",
   178 => x"80c6d00c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b0bbf",
   183 => x"900c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80c6d0",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80c6",
   208 => x"b80c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050d84bf",
   216 => x"5186c72d",
   217 => x"ff115170",
   218 => x"8025f638",
   219 => x"0284050d",
   220 => x"0402fc05",
   221 => x"0dec5183",
   222 => x"710c86c7",
   223 => x"2d82710c",
   224 => x"90a42d02",
   225 => x"84050d04",
   226 => x"02fc050d",
   227 => x"ec518182",
   228 => x"710c86c7",
   229 => x"2d82710c",
   230 => x"90a42d02",
   231 => x"84050d04",
   232 => x"02fc050d",
   233 => x"ec5180c2",
   234 => x"710c86c7",
   235 => x"2d82710c",
   236 => x"90a42d02",
   237 => x"84050d04",
   238 => x"02fc050d",
   239 => x"ec518282",
   240 => x"710c86c7",
   241 => x"2d82710c",
   242 => x"90a42d02",
   243 => x"84050d04",
   244 => x"02fc050d",
   245 => x"ec519271",
   246 => x"0c86c72d",
   247 => x"82710c02",
   248 => x"84050d04",
   249 => x"02d0050d",
   250 => x"7d548074",
   251 => x"5380c6d4",
   252 => x"525bab8a",
   253 => x"2d80c6b8",
   254 => x"087b2e81",
   255 => x"b63880c6",
   256 => x"d80870f8",
   257 => x"0c891580",
   258 => x"f52d8a16",
   259 => x"80f52d71",
   260 => x"82802905",
   261 => x"881780f5",
   262 => x"2d708480",
   263 => x"802912f4",
   264 => x"0c575556",
   265 => x"58a40bec",
   266 => x"0c7aff19",
   267 => x"585a767b",
   268 => x"2e8b3881",
   269 => x"1a77812a",
   270 => x"585a76f7",
   271 => x"38f71a5a",
   272 => x"815b8078",
   273 => x"2580ec38",
   274 => x"79527651",
   275 => x"84a82d80",
   276 => x"c7a05280",
   277 => x"c6d451ad",
   278 => x"d72d80c6",
   279 => x"b808802e",
   280 => x"b93880c7",
   281 => x"a05c83fc",
   282 => x"597b7084",
   283 => x"055d0870",
   284 => x"81ff0671",
   285 => x"882a7081",
   286 => x"ff067390",
   287 => x"2a7081ff",
   288 => x"0675982a",
   289 => x"e80ce80c",
   290 => x"58e80c57",
   291 => x"e80cfc1a",
   292 => x"5a537880",
   293 => x"25d33889",
   294 => x"a20480c6",
   295 => x"b8085b84",
   296 => x"805880c6",
   297 => x"d451ada7",
   298 => x"2dfc8018",
   299 => x"81185858",
   300 => x"88c20486",
   301 => x"da2d840b",
   302 => x"ec0c7a80",
   303 => x"2e8e3880",
   304 => x"c2a85192",
   305 => x"ae2d90a4",
   306 => x"2d89d304",
   307 => x"80c48851",
   308 => x"92ae2d7a",
   309 => x"80c6b80c",
   310 => x"02b0050d",
   311 => x"0402ec05",
   312 => x"0d840bec",
   313 => x"0c90822d",
   314 => x"8cd42d81",
   315 => x"f92da1ca",
   316 => x"2d80c6b8",
   317 => x"08802e82",
   318 => x"c43887e4",
   319 => x"51b4972d",
   320 => x"80c2a851",
   321 => x"92ae2d90",
   322 => x"a42d8ce0",
   323 => x"2d92c12d",
   324 => x"80c1b00b",
   325 => x"80f52d70",
   326 => x"822b8406",
   327 => x"80c1bc0b",
   328 => x"80f52d70",
   329 => x"982b8180",
   330 => x"0a0680c1",
   331 => x"c80b80f5",
   332 => x"2d70842b",
   333 => x"b0067473",
   334 => x"070780c1",
   335 => x"d40b80f5",
   336 => x"2d70882b",
   337 => x"8e800680",
   338 => x"c08c0b80",
   339 => x"f52d708d",
   340 => x"2b80c080",
   341 => x"06747307",
   342 => x"0780c098",
   343 => x"0b80f52d",
   344 => x"70902b84",
   345 => x"80800680",
   346 => x"c0a40b80",
   347 => x"f52d7094",
   348 => x"2b9c800a",
   349 => x"06747307",
   350 => x"0780c0b0",
   351 => x"0b80f52d",
   352 => x"70862b80",
   353 => x"c00680c0",
   354 => x"bc0b80f5",
   355 => x"2d708c2b",
   356 => x"a0800674",
   357 => x"73070780",
   358 => x"c0c80b80",
   359 => x"f52d7092",
   360 => x"2bb08080",
   361 => x"06bf9c0b",
   362 => x"80f52d70",
   363 => x"832b8806",
   364 => x"74730707",
   365 => x"bfa80b80",
   366 => x"f52d7010",
   367 => x"8206bfb4",
   368 => x"0b80f52d",
   369 => x"709a2bb0",
   370 => x"0a067473",
   371 => x"0707bfc0",
   372 => x"0b80f52d",
   373 => x"709c2b8c",
   374 => x"0a0680c3",
   375 => x"900b80f5",
   376 => x"2d708e2b",
   377 => x"83808006",
   378 => x"74730707",
   379 => x"80c39c0b",
   380 => x"80f52d70",
   381 => x"8b2b9080",
   382 => x"0680c3a8",
   383 => x"0b80f52d",
   384 => x"709e2b82",
   385 => x"0a067473",
   386 => x"0707fc0c",
   387 => x"54545454",
   388 => x"54545454",
   389 => x"54545454",
   390 => x"54545454",
   391 => x"54545454",
   392 => x"54545454",
   393 => x"54545654",
   394 => x"52575753",
   395 => x"53865280",
   396 => x"c6b80883",
   397 => x"38845271",
   398 => x"ec0c8a8a",
   399 => x"04800b80",
   400 => x"c6b80c02",
   401 => x"94050d04",
   402 => x"71980c04",
   403 => x"ffb00880",
   404 => x"c6b80c04",
   405 => x"810bffb0",
   406 => x"0c04800b",
   407 => x"ffb00c04",
   408 => x"02f4050d",
   409 => x"8dee0480",
   410 => x"c6b80881",
   411 => x"f02e0981",
   412 => x"068a3881",
   413 => x"0b80c4ec",
   414 => x"0c8dee04",
   415 => x"80c6b808",
   416 => x"81e02e09",
   417 => x"81068a38",
   418 => x"810b80c4",
   419 => x"f00c8dee",
   420 => x"0480c6b8",
   421 => x"085280c4",
   422 => x"f008802e",
   423 => x"893880c6",
   424 => x"b8088180",
   425 => x"05527184",
   426 => x"2c728f06",
   427 => x"535380c4",
   428 => x"ec08802e",
   429 => x"9a387284",
   430 => x"2980c4ac",
   431 => x"05721381",
   432 => x"712b7009",
   433 => x"73080673",
   434 => x"0c515353",
   435 => x"8de20472",
   436 => x"842980c4",
   437 => x"ac057213",
   438 => x"83712b72",
   439 => x"0807720c",
   440 => x"5353800b",
   441 => x"80c4f00c",
   442 => x"800b80c4",
   443 => x"ec0c80c6",
   444 => x"e0518ef5",
   445 => x"2d80c6b8",
   446 => x"08ff24fe",
   447 => x"ea38800b",
   448 => x"80c6b80c",
   449 => x"028c050d",
   450 => x"0402f805",
   451 => x"0d80c4ac",
   452 => x"528f5180",
   453 => x"72708405",
   454 => x"540cff11",
   455 => x"51708025",
   456 => x"f2380288",
   457 => x"050d0402",
   458 => x"f0050d75",
   459 => x"518cda2d",
   460 => x"70822cfc",
   461 => x"0680c4ac",
   462 => x"1172109e",
   463 => x"06710870",
   464 => x"722a7083",
   465 => x"0682742b",
   466 => x"70097406",
   467 => x"760c5451",
   468 => x"56575351",
   469 => x"538cd42d",
   470 => x"7180c6b8",
   471 => x"0c029005",
   472 => x"0d0402fc",
   473 => x"050d7251",
   474 => x"80710c80",
   475 => x"0b84120c",
   476 => x"0284050d",
   477 => x"0402f005",
   478 => x"0d757008",
   479 => x"84120853",
   480 => x"5353ff54",
   481 => x"71712ea8",
   482 => x"388cda2d",
   483 => x"84130870",
   484 => x"84291488",
   485 => x"11700870",
   486 => x"81ff0684",
   487 => x"18088111",
   488 => x"8706841a",
   489 => x"0c535155",
   490 => x"5151518c",
   491 => x"d42d7154",
   492 => x"7380c6b8",
   493 => x"0c029005",
   494 => x"0d0402f8",
   495 => x"050d8cda",
   496 => x"2de00870",
   497 => x"8b2a7081",
   498 => x"06515252",
   499 => x"70802ea1",
   500 => x"3880c6e0",
   501 => x"08708429",
   502 => x"80c6e805",
   503 => x"7381ff06",
   504 => x"710c5151",
   505 => x"80c6e008",
   506 => x"81118706",
   507 => x"80c6e00c",
   508 => x"51800b80",
   509 => x"c7880c8c",
   510 => x"cc2d8cd4",
   511 => x"2d028805",
   512 => x"0d0402fc",
   513 => x"050d80c6",
   514 => x"e0518ee2",
   515 => x"2d8e892d",
   516 => x"8fba518c",
   517 => x"c82d0284",
   518 => x"050d0480",
   519 => x"c78c0880",
   520 => x"c6b80c04",
   521 => x"02fc050d",
   522 => x"90ae048c",
   523 => x"e02d80f6",
   524 => x"518ea72d",
   525 => x"80c6b808",
   526 => x"f23880da",
   527 => x"518ea72d",
   528 => x"80c6b808",
   529 => x"e63880c6",
   530 => x"b80880c4",
   531 => x"f80c80c6",
   532 => x"b8085185",
   533 => x"8d2d0284",
   534 => x"050d0402",
   535 => x"ec050d76",
   536 => x"54805287",
   537 => x"0b881580",
   538 => x"f52d5653",
   539 => x"74722483",
   540 => x"38a05372",
   541 => x"5183842d",
   542 => x"81128b15",
   543 => x"80f52d54",
   544 => x"52727225",
   545 => x"de380294",
   546 => x"050d0402",
   547 => x"f0050d80",
   548 => x"c78c0854",
   549 => x"81f92d80",
   550 => x"0b80c790",
   551 => x"0c730880",
   552 => x"2e818638",
   553 => x"820b80c6",
   554 => x"cc0c80c7",
   555 => x"90088f06",
   556 => x"80c6c80c",
   557 => x"73085271",
   558 => x"832e9638",
   559 => x"71832689",
   560 => x"3871812e",
   561 => x"af389292",
   562 => x"0471852e",
   563 => x"9f389292",
   564 => x"04881480",
   565 => x"f52d8415",
   566 => x"08bddc53",
   567 => x"545286a0",
   568 => x"2d718429",
   569 => x"13700852",
   570 => x"52929604",
   571 => x"735190db",
   572 => x"2d929204",
   573 => x"80c4f408",
   574 => x"8815082c",
   575 => x"70810651",
   576 => x"5271802e",
   577 => x"8738bde0",
   578 => x"51928f04",
   579 => x"bde45186",
   580 => x"a02d8414",
   581 => x"085186a0",
   582 => x"2d80c790",
   583 => x"08810580",
   584 => x"c7900c8c",
   585 => x"1454919d",
   586 => x"04029005",
   587 => x"0d047180",
   588 => x"c78c0c91",
   589 => x"8b2d80c7",
   590 => x"9008ff05",
   591 => x"80c7940c",
   592 => x"0402e805",
   593 => x"0d80c78c",
   594 => x"0880c798",
   595 => x"08575587",
   596 => x"518ea72d",
   597 => x"80c6b808",
   598 => x"812a7081",
   599 => x"06515271",
   600 => x"802ea338",
   601 => x"92ea048c",
   602 => x"e02d8751",
   603 => x"8ea72d80",
   604 => x"c6b808f3",
   605 => x"3880c4f8",
   606 => x"08813270",
   607 => x"80c4f80c",
   608 => x"70525285",
   609 => x"8d2d80fe",
   610 => x"518ea72d",
   611 => x"80c6b808",
   612 => x"802ea938",
   613 => x"80c4f808",
   614 => x"802e9238",
   615 => x"800b80c4",
   616 => x"f80c8051",
   617 => x"858d2d93",
   618 => x"ad048ce0",
   619 => x"2d80fe51",
   620 => x"8ea72d80",
   621 => x"c6b808f2",
   622 => x"3887d02d",
   623 => x"80c4f808",
   624 => x"903881fd",
   625 => x"518ea72d",
   626 => x"81fa518e",
   627 => x"a72d99a6",
   628 => x"0481f551",
   629 => x"8ea72d80",
   630 => x"c6b80881",
   631 => x"2a708106",
   632 => x"51527180",
   633 => x"2eb33880",
   634 => x"c7940852",
   635 => x"71802e8a",
   636 => x"38ff1280",
   637 => x"c7940c94",
   638 => x"990480c7",
   639 => x"90081080",
   640 => x"c7900805",
   641 => x"70842916",
   642 => x"51528812",
   643 => x"08802e89",
   644 => x"38ff5188",
   645 => x"12085271",
   646 => x"2d81f251",
   647 => x"8ea72d80",
   648 => x"c6b80881",
   649 => x"2a708106",
   650 => x"51527180",
   651 => x"2eb43880",
   652 => x"c79008ff",
   653 => x"1180c794",
   654 => x"08565353",
   655 => x"7372258a",
   656 => x"38811480",
   657 => x"c7940c94",
   658 => x"e2047210",
   659 => x"13708429",
   660 => x"16515288",
   661 => x"1208802e",
   662 => x"8938fe51",
   663 => x"88120852",
   664 => x"712d81fd",
   665 => x"518ea72d",
   666 => x"80c6b808",
   667 => x"812a7081",
   668 => x"06515271",
   669 => x"802eb138",
   670 => x"80c79408",
   671 => x"802e8a38",
   672 => x"800b80c7",
   673 => x"940c95a8",
   674 => x"0480c790",
   675 => x"081080c7",
   676 => x"90080570",
   677 => x"84291651",
   678 => x"52881208",
   679 => x"802e8938",
   680 => x"fd518812",
   681 => x"0852712d",
   682 => x"81fa518e",
   683 => x"a72d80c6",
   684 => x"b808812a",
   685 => x"70810651",
   686 => x"5271802e",
   687 => x"b13880c7",
   688 => x"9008ff11",
   689 => x"545280c7",
   690 => x"94087325",
   691 => x"89387280",
   692 => x"c7940c95",
   693 => x"ee047110",
   694 => x"12708429",
   695 => x"16515288",
   696 => x"1208802e",
   697 => x"8938fc51",
   698 => x"88120852",
   699 => x"712d80c7",
   700 => x"94087053",
   701 => x"5473802e",
   702 => x"8a388c15",
   703 => x"ff155555",
   704 => x"95f50482",
   705 => x"0b80c6cc",
   706 => x"0c718f06",
   707 => x"80c6c80c",
   708 => x"81eb518e",
   709 => x"a72d80c6",
   710 => x"b808812a",
   711 => x"70810651",
   712 => x"5271802e",
   713 => x"ad387408",
   714 => x"852e0981",
   715 => x"06a43888",
   716 => x"1580f52d",
   717 => x"ff055271",
   718 => x"881681b7",
   719 => x"2d71982b",
   720 => x"52718025",
   721 => x"8838800b",
   722 => x"881681b7",
   723 => x"2d745190",
   724 => x"db2d81f4",
   725 => x"518ea72d",
   726 => x"80c6b808",
   727 => x"812a7081",
   728 => x"06515271",
   729 => x"802eb338",
   730 => x"7408852e",
   731 => x"098106aa",
   732 => x"38881580",
   733 => x"f52d8105",
   734 => x"52718816",
   735 => x"81b72d71",
   736 => x"81ff068b",
   737 => x"1680f52d",
   738 => x"54527272",
   739 => x"27873872",
   740 => x"881681b7",
   741 => x"2d745190",
   742 => x"db2d80da",
   743 => x"518ea72d",
   744 => x"80c6b808",
   745 => x"812a7081",
   746 => x"06515271",
   747 => x"802e81ad",
   748 => x"3880c78c",
   749 => x"0880c794",
   750 => x"08555373",
   751 => x"802e8a38",
   752 => x"8c13ff15",
   753 => x"555397bb",
   754 => x"04720852",
   755 => x"71822ea6",
   756 => x"38718226",
   757 => x"89387181",
   758 => x"2eaa3898",
   759 => x"dd047183",
   760 => x"2eb43871",
   761 => x"842e0981",
   762 => x"0680f238",
   763 => x"88130851",
   764 => x"92ae2d98",
   765 => x"dd0480c7",
   766 => x"94085188",
   767 => x"13085271",
   768 => x"2d98dd04",
   769 => x"810b8814",
   770 => x"082b80c4",
   771 => x"f4083280",
   772 => x"c4f40c98",
   773 => x"b1048813",
   774 => x"80f52d81",
   775 => x"058b1480",
   776 => x"f52d5354",
   777 => x"71742483",
   778 => x"38805473",
   779 => x"881481b7",
   780 => x"2d918b2d",
   781 => x"98dd0475",
   782 => x"08802ea4",
   783 => x"38750851",
   784 => x"8ea72d80",
   785 => x"c6b80881",
   786 => x"06527180",
   787 => x"2e8c3880",
   788 => x"c7940851",
   789 => x"84160852",
   790 => x"712d8816",
   791 => x"5675d838",
   792 => x"8054800b",
   793 => x"80c6cc0c",
   794 => x"738f0680",
   795 => x"c6c80ca0",
   796 => x"527380c7",
   797 => x"94082e09",
   798 => x"81069938",
   799 => x"80c79008",
   800 => x"ff057432",
   801 => x"70098105",
   802 => x"7072079f",
   803 => x"2a917131",
   804 => x"51515353",
   805 => x"71518384",
   806 => x"2d811454",
   807 => x"8e7425c2",
   808 => x"3880c4f8",
   809 => x"08527180",
   810 => x"c6b80c02",
   811 => x"98050d04",
   812 => x"02f4050d",
   813 => x"d45281ff",
   814 => x"720c7108",
   815 => x"5381ff72",
   816 => x"0c72882b",
   817 => x"83fe8006",
   818 => x"72087081",
   819 => x"ff065152",
   820 => x"5381ff72",
   821 => x"0c727107",
   822 => x"882b7208",
   823 => x"7081ff06",
   824 => x"51525381",
   825 => x"ff720c72",
   826 => x"7107882b",
   827 => x"72087081",
   828 => x"ff067207",
   829 => x"80c6b80c",
   830 => x"5253028c",
   831 => x"050d0402",
   832 => x"f4050d74",
   833 => x"767181ff",
   834 => x"06d40c53",
   835 => x"5380c79c",
   836 => x"08853871",
   837 => x"892b5271",
   838 => x"982ad40c",
   839 => x"71902a70",
   840 => x"81ff06d4",
   841 => x"0c517188",
   842 => x"2a7081ff",
   843 => x"06d40c51",
   844 => x"7181ff06",
   845 => x"d40c7290",
   846 => x"2a7081ff",
   847 => x"06d40c51",
   848 => x"d4087081",
   849 => x"ff065151",
   850 => x"82b8bf52",
   851 => x"7081ff2e",
   852 => x"09810694",
   853 => x"3881ff0b",
   854 => x"d40cd408",
   855 => x"7081ff06",
   856 => x"ff145451",
   857 => x"5171e538",
   858 => x"7080c6b8",
   859 => x"0c028c05",
   860 => x"0d0402fc",
   861 => x"050d81c7",
   862 => x"5181ff0b",
   863 => x"d40cff11",
   864 => x"51708025",
   865 => x"f4380284",
   866 => x"050d0402",
   867 => x"f4050d81",
   868 => x"ff0bd40c",
   869 => x"93538052",
   870 => x"87fc80c1",
   871 => x"5199ff2d",
   872 => x"80c6b808",
   873 => x"8b3881ff",
   874 => x"0bd40c81",
   875 => x"539bb904",
   876 => x"9af22dff",
   877 => x"135372de",
   878 => x"387280c6",
   879 => x"b80c028c",
   880 => x"050d0402",
   881 => x"ec050d81",
   882 => x"0b80c79c",
   883 => x"0c8454d0",
   884 => x"08708f2a",
   885 => x"70810651",
   886 => x"515372f3",
   887 => x"3872d00c",
   888 => x"9af22dbd",
   889 => x"e85186a0",
   890 => x"2dd00870",
   891 => x"8f2a7081",
   892 => x"06515153",
   893 => x"72f33881",
   894 => x"0bd00cb1",
   895 => x"53805284",
   896 => x"d480c051",
   897 => x"99ff2d80",
   898 => x"c6b80881",
   899 => x"2e933872",
   900 => x"822ebf38",
   901 => x"ff135372",
   902 => x"e438ff14",
   903 => x"5473ffaf",
   904 => x"389af22d",
   905 => x"83aa5284",
   906 => x"9c80c851",
   907 => x"99ff2d80",
   908 => x"c6b80881",
   909 => x"2e098106",
   910 => x"933899b0",
   911 => x"2d80c6b8",
   912 => x"0883ffff",
   913 => x"06537283",
   914 => x"aa2e9d38",
   915 => x"9b8b2d9c",
   916 => x"e304bdf4",
   917 => x"5186a02d",
   918 => x"80539eb8",
   919 => x"04be8c51",
   920 => x"86a02d80",
   921 => x"549e8904",
   922 => x"81ff0bd4",
   923 => x"0cb1549a",
   924 => x"f22d8fcf",
   925 => x"53805287",
   926 => x"fc80f751",
   927 => x"99ff2d80",
   928 => x"c6b80855",
   929 => x"80c6b808",
   930 => x"812e0981",
   931 => x"069c3881",
   932 => x"ff0bd40c",
   933 => x"820a5284",
   934 => x"9c80e951",
   935 => x"99ff2d80",
   936 => x"c6b80880",
   937 => x"2e8d389a",
   938 => x"f22dff13",
   939 => x"5372c638",
   940 => x"9dfc0481",
   941 => x"ff0bd40c",
   942 => x"80c6b808",
   943 => x"5287fc80",
   944 => x"fa5199ff",
   945 => x"2d80c6b8",
   946 => x"08b23881",
   947 => x"ff0bd40c",
   948 => x"d4085381",
   949 => x"ff0bd40c",
   950 => x"81ff0bd4",
   951 => x"0c81ff0b",
   952 => x"d40c81ff",
   953 => x"0bd40c72",
   954 => x"862a7081",
   955 => x"06765651",
   956 => x"53729638",
   957 => x"80c6b808",
   958 => x"549e8904",
   959 => x"73822efe",
   960 => x"dc38ff14",
   961 => x"5473fee7",
   962 => x"387380c7",
   963 => x"9c0c738b",
   964 => x"38815287",
   965 => x"fc80d051",
   966 => x"99ff2d81",
   967 => x"ff0bd40c",
   968 => x"d008708f",
   969 => x"2a708106",
   970 => x"51515372",
   971 => x"f33872d0",
   972 => x"0c81ff0b",
   973 => x"d40c8153",
   974 => x"7280c6b8",
   975 => x"0c029405",
   976 => x"0d0402e8",
   977 => x"050d7855",
   978 => x"805681ff",
   979 => x"0bd40cd0",
   980 => x"08708f2a",
   981 => x"70810651",
   982 => x"515372f3",
   983 => x"3882810b",
   984 => x"d00c81ff",
   985 => x"0bd40c77",
   986 => x"5287fc80",
   987 => x"d15199ff",
   988 => x"2d80dbc6",
   989 => x"df5480c6",
   990 => x"b808802e",
   991 => x"8a38beac",
   992 => x"5186a02d",
   993 => x"9fdb0481",
   994 => x"ff0bd40c",
   995 => x"d4087081",
   996 => x"ff065153",
   997 => x"7281fe2e",
   998 => x"0981069e",
   999 => x"3880ff53",
  1000 => x"99b02d80",
  1001 => x"c6b80875",
  1002 => x"70840557",
  1003 => x"0cff1353",
  1004 => x"728025ec",
  1005 => x"3881569f",
  1006 => x"c004ff14",
  1007 => x"5473c838",
  1008 => x"81ff0bd4",
  1009 => x"0c81ff0b",
  1010 => x"d40cd008",
  1011 => x"708f2a70",
  1012 => x"81065151",
  1013 => x"5372f338",
  1014 => x"72d00c75",
  1015 => x"80c6b80c",
  1016 => x"0298050d",
  1017 => x"0402e805",
  1018 => x"0d77797b",
  1019 => x"58555580",
  1020 => x"53727625",
  1021 => x"a3387470",
  1022 => x"81055680",
  1023 => x"f52d7470",
  1024 => x"81055680",
  1025 => x"f52d5252",
  1026 => x"71712e86",
  1027 => x"388151a0",
  1028 => x"9a048113",
  1029 => x"539ff104",
  1030 => x"80517080",
  1031 => x"c6b80c02",
  1032 => x"98050d04",
  1033 => x"02ec050d",
  1034 => x"76557480",
  1035 => x"2e80c238",
  1036 => x"9a1580e0",
  1037 => x"2d51aeb1",
  1038 => x"2d80c6b8",
  1039 => x"0880c6b8",
  1040 => x"0880cdd0",
  1041 => x"0c80c6b8",
  1042 => x"08545480",
  1043 => x"cdac0880",
  1044 => x"2e9a3894",
  1045 => x"1580e02d",
  1046 => x"51aeb12d",
  1047 => x"80c6b808",
  1048 => x"902b83ff",
  1049 => x"f00a0670",
  1050 => x"75075153",
  1051 => x"7280cdd0",
  1052 => x"0c80cdd0",
  1053 => x"08537280",
  1054 => x"2e9d3880",
  1055 => x"cda408fe",
  1056 => x"14712980",
  1057 => x"cdb80805",
  1058 => x"80cdd40c",
  1059 => x"70842b80",
  1060 => x"cdb00c54",
  1061 => x"a1c50480",
  1062 => x"cdbc0880",
  1063 => x"cdd00c80",
  1064 => x"cdc00880",
  1065 => x"cdd40c80",
  1066 => x"cdac0880",
  1067 => x"2e8b3880",
  1068 => x"cda40884",
  1069 => x"2b53a1c0",
  1070 => x"0480cdc4",
  1071 => x"08842b53",
  1072 => x"7280cdb0",
  1073 => x"0c029405",
  1074 => x"0d0402d8",
  1075 => x"050d800b",
  1076 => x"80cdac0c",
  1077 => x"84549bc3",
  1078 => x"2d80c6b8",
  1079 => x"08802e97",
  1080 => x"3880c7a0",
  1081 => x"5280519e",
  1082 => x"c22d80c6",
  1083 => x"b808802e",
  1084 => x"8638fe54",
  1085 => x"a1ff04ff",
  1086 => x"14547380",
  1087 => x"24d83873",
  1088 => x"8c38bebc",
  1089 => x"5186a02d",
  1090 => x"7355a7cc",
  1091 => x"04805681",
  1092 => x"0b80cdd8",
  1093 => x"0c8853be",
  1094 => x"d05280c7",
  1095 => x"d6519fe5",
  1096 => x"2d80c6b8",
  1097 => x"08762e09",
  1098 => x"81068938",
  1099 => x"80c6b808",
  1100 => x"80cdd80c",
  1101 => x"8853bedc",
  1102 => x"5280c7f2",
  1103 => x"519fe52d",
  1104 => x"80c6b808",
  1105 => x"893880c6",
  1106 => x"b80880cd",
  1107 => x"d80c80cd",
  1108 => x"d808802e",
  1109 => x"81803880",
  1110 => x"cae60b80",
  1111 => x"f52d80ca",
  1112 => x"e70b80f5",
  1113 => x"2d71982b",
  1114 => x"71902b07",
  1115 => x"80cae80b",
  1116 => x"80f52d70",
  1117 => x"882b7207",
  1118 => x"80cae90b",
  1119 => x"80f52d71",
  1120 => x"0780cb9e",
  1121 => x"0b80f52d",
  1122 => x"80cb9f0b",
  1123 => x"80f52d71",
  1124 => x"882b0753",
  1125 => x"5f54525a",
  1126 => x"56575573",
  1127 => x"81abaa2e",
  1128 => x"0981068e",
  1129 => x"387551ae",
  1130 => x"802d80c6",
  1131 => x"b80856a3",
  1132 => x"bf047382",
  1133 => x"d4d52e87",
  1134 => x"38bee851",
  1135 => x"a4880480",
  1136 => x"c7a05275",
  1137 => x"519ec22d",
  1138 => x"80c6b808",
  1139 => x"5580c6b8",
  1140 => x"08802e83",
  1141 => x"f7388853",
  1142 => x"bedc5280",
  1143 => x"c7f2519f",
  1144 => x"e52d80c6",
  1145 => x"b8088a38",
  1146 => x"810b80cd",
  1147 => x"ac0ca48e",
  1148 => x"048853be",
  1149 => x"d05280c7",
  1150 => x"d6519fe5",
  1151 => x"2d80c6b8",
  1152 => x"08802e8a",
  1153 => x"38befc51",
  1154 => x"86a02da4",
  1155 => x"ed0480cb",
  1156 => x"9e0b80f5",
  1157 => x"2d547380",
  1158 => x"d52e0981",
  1159 => x"0680ce38",
  1160 => x"80cb9f0b",
  1161 => x"80f52d54",
  1162 => x"7381aa2e",
  1163 => x"098106bd",
  1164 => x"38800b80",
  1165 => x"c7a00b80",
  1166 => x"f52d5654",
  1167 => x"7481e92e",
  1168 => x"83388154",
  1169 => x"7481eb2e",
  1170 => x"8c388055",
  1171 => x"73752e09",
  1172 => x"810682f8",
  1173 => x"3880c7ab",
  1174 => x"0b80f52d",
  1175 => x"55748e38",
  1176 => x"80c7ac0b",
  1177 => x"80f52d54",
  1178 => x"73822e86",
  1179 => x"388055a7",
  1180 => x"cc0480c7",
  1181 => x"ad0b80f5",
  1182 => x"2d7080cd",
  1183 => x"a40cff05",
  1184 => x"80cda80c",
  1185 => x"80c7ae0b",
  1186 => x"80f52d80",
  1187 => x"c7af0b80",
  1188 => x"f52d5876",
  1189 => x"05778280",
  1190 => x"29057080",
  1191 => x"cdb40c80",
  1192 => x"c7b00b80",
  1193 => x"f52d7080",
  1194 => x"cdc80c80",
  1195 => x"cdac0859",
  1196 => x"57587680",
  1197 => x"2e81b638",
  1198 => x"8853bedc",
  1199 => x"5280c7f2",
  1200 => x"519fe52d",
  1201 => x"80c6b808",
  1202 => x"82823880",
  1203 => x"cda40870",
  1204 => x"842b80cd",
  1205 => x"b00c7080",
  1206 => x"cdc40c80",
  1207 => x"c7c50b80",
  1208 => x"f52d80c7",
  1209 => x"c40b80f5",
  1210 => x"2d718280",
  1211 => x"290580c7",
  1212 => x"c60b80f5",
  1213 => x"2d708480",
  1214 => x"80291280",
  1215 => x"c7c70b80",
  1216 => x"f52d7081",
  1217 => x"800a2912",
  1218 => x"7080cdcc",
  1219 => x"0c80cdc8",
  1220 => x"08712980",
  1221 => x"cdb40805",
  1222 => x"7080cdb8",
  1223 => x"0c80c7cd",
  1224 => x"0b80f52d",
  1225 => x"80c7cc0b",
  1226 => x"80f52d71",
  1227 => x"82802905",
  1228 => x"80c7ce0b",
  1229 => x"80f52d70",
  1230 => x"84808029",
  1231 => x"1280c7cf",
  1232 => x"0b80f52d",
  1233 => x"70982b81",
  1234 => x"f00a0672",
  1235 => x"057080cd",
  1236 => x"bc0cfe11",
  1237 => x"7e297705",
  1238 => x"80cdc00c",
  1239 => x"52595243",
  1240 => x"545e5152",
  1241 => x"59525d57",
  1242 => x"5957a7c5",
  1243 => x"0480c7b2",
  1244 => x"0b80f52d",
  1245 => x"80c7b10b",
  1246 => x"80f52d71",
  1247 => x"82802905",
  1248 => x"7080cdb0",
  1249 => x"0c70a029",
  1250 => x"83ff0570",
  1251 => x"892a7080",
  1252 => x"cdc40c80",
  1253 => x"c7b70b80",
  1254 => x"f52d80c7",
  1255 => x"b60b80f5",
  1256 => x"2d718280",
  1257 => x"29057080",
  1258 => x"cdcc0c7b",
  1259 => x"71291e70",
  1260 => x"80cdc00c",
  1261 => x"7d80cdbc",
  1262 => x"0c730580",
  1263 => x"cdb80c55",
  1264 => x"5e515155",
  1265 => x"558051a0",
  1266 => x"a42d8155",
  1267 => x"7480c6b8",
  1268 => x"0c02a805",
  1269 => x"0d0402ec",
  1270 => x"050d7670",
  1271 => x"872c7180",
  1272 => x"ff065556",
  1273 => x"5480cdac",
  1274 => x"088a3873",
  1275 => x"882c7481",
  1276 => x"ff065455",
  1277 => x"80c7a052",
  1278 => x"80cdb408",
  1279 => x"15519ec2",
  1280 => x"2d80c6b8",
  1281 => x"085480c6",
  1282 => x"b808802e",
  1283 => x"b83880cd",
  1284 => x"ac08802e",
  1285 => x"9a387284",
  1286 => x"2980c7a0",
  1287 => x"05700852",
  1288 => x"53ae802d",
  1289 => x"80c6b808",
  1290 => x"f00a0653",
  1291 => x"a8c30472",
  1292 => x"1080c7a0",
  1293 => x"057080e0",
  1294 => x"2d5253ae",
  1295 => x"b12d80c6",
  1296 => x"b8085372",
  1297 => x"547380c6",
  1298 => x"b80c0294",
  1299 => x"050d0402",
  1300 => x"e0050d79",
  1301 => x"70842c80",
  1302 => x"cdd40805",
  1303 => x"718f0652",
  1304 => x"5553728a",
  1305 => x"3880c7a0",
  1306 => x"5273519e",
  1307 => x"c22d72a0",
  1308 => x"2980c7a0",
  1309 => x"05548074",
  1310 => x"80f52d56",
  1311 => x"5374732e",
  1312 => x"83388153",
  1313 => x"7481e52e",
  1314 => x"81f43881",
  1315 => x"70740654",
  1316 => x"5872802e",
  1317 => x"81e8388b",
  1318 => x"1480f52d",
  1319 => x"70832a79",
  1320 => x"06585676",
  1321 => x"9b3880c4",
  1322 => x"fc085372",
  1323 => x"89387280",
  1324 => x"cba00b81",
  1325 => x"b72d7680",
  1326 => x"c4fc0c73",
  1327 => x"53ab8004",
  1328 => x"758f2e09",
  1329 => x"810681b6",
  1330 => x"38749f06",
  1331 => x"8d2980cb",
  1332 => x"93115153",
  1333 => x"811480f5",
  1334 => x"2d737081",
  1335 => x"055581b7",
  1336 => x"2d831480",
  1337 => x"f52d7370",
  1338 => x"81055581",
  1339 => x"b72d8514",
  1340 => x"80f52d73",
  1341 => x"70810555",
  1342 => x"81b72d87",
  1343 => x"1480f52d",
  1344 => x"73708105",
  1345 => x"5581b72d",
  1346 => x"891480f5",
  1347 => x"2d737081",
  1348 => x"055581b7",
  1349 => x"2d8e1480",
  1350 => x"f52d7370",
  1351 => x"81055581",
  1352 => x"b72d9014",
  1353 => x"80f52d73",
  1354 => x"70810555",
  1355 => x"81b72d92",
  1356 => x"1480f52d",
  1357 => x"73708105",
  1358 => x"5581b72d",
  1359 => x"941480f5",
  1360 => x"2d737081",
  1361 => x"055581b7",
  1362 => x"2d961480",
  1363 => x"f52d7370",
  1364 => x"81055581",
  1365 => x"b72d9814",
  1366 => x"80f52d73",
  1367 => x"70810555",
  1368 => x"81b72d9c",
  1369 => x"1480f52d",
  1370 => x"73708105",
  1371 => x"5581b72d",
  1372 => x"9e1480f5",
  1373 => x"2d7381b7",
  1374 => x"2d7780c4",
  1375 => x"fc0c8053",
  1376 => x"7280c6b8",
  1377 => x"0c02a005",
  1378 => x"0d0402cc",
  1379 => x"050d7e60",
  1380 => x"5e5a800b",
  1381 => x"80cdd008",
  1382 => x"80cdd408",
  1383 => x"595c5680",
  1384 => x"5880cdb0",
  1385 => x"08782e81",
  1386 => x"b838778f",
  1387 => x"06a01757",
  1388 => x"54739138",
  1389 => x"80c7a052",
  1390 => x"76518117",
  1391 => x"579ec22d",
  1392 => x"80c7a056",
  1393 => x"807680f5",
  1394 => x"2d565474",
  1395 => x"742e8338",
  1396 => x"81547481",
  1397 => x"e52e80fd",
  1398 => x"38817075",
  1399 => x"06555c73",
  1400 => x"802e80f1",
  1401 => x"388b1680",
  1402 => x"f52d9806",
  1403 => x"597880e5",
  1404 => x"388b537c",
  1405 => x"5275519f",
  1406 => x"e52d80c6",
  1407 => x"b80880d5",
  1408 => x"389c1608",
  1409 => x"51ae802d",
  1410 => x"80c6b808",
  1411 => x"841b0c9a",
  1412 => x"1680e02d",
  1413 => x"51aeb12d",
  1414 => x"80c6b808",
  1415 => x"80c6b808",
  1416 => x"881c0c80",
  1417 => x"c6b80855",
  1418 => x"5580cdac",
  1419 => x"08802e99",
  1420 => x"38941680",
  1421 => x"e02d51ae",
  1422 => x"b12d80c6",
  1423 => x"b808902b",
  1424 => x"83fff00a",
  1425 => x"06701651",
  1426 => x"5473881b",
  1427 => x"0c787a0c",
  1428 => x"7b54ad9d",
  1429 => x"04811858",
  1430 => x"80cdb008",
  1431 => x"7826feca",
  1432 => x"3880cdac",
  1433 => x"08802eb3",
  1434 => x"387a51a7",
  1435 => x"d62d80c6",
  1436 => x"b80880c6",
  1437 => x"b80880ff",
  1438 => x"fffff806",
  1439 => x"555b7380",
  1440 => x"fffffff8",
  1441 => x"2e953880",
  1442 => x"c6b808fe",
  1443 => x"0580cda4",
  1444 => x"082980cd",
  1445 => x"b8080557",
  1446 => x"ab9f0480",
  1447 => x"547380c6",
  1448 => x"b80c02b4",
  1449 => x"050d0402",
  1450 => x"f4050d74",
  1451 => x"70088105",
  1452 => x"710c7008",
  1453 => x"80cda808",
  1454 => x"06535371",
  1455 => x"8f388813",
  1456 => x"0851a7d6",
  1457 => x"2d80c6b8",
  1458 => x"0888140c",
  1459 => x"810b80c6",
  1460 => x"b80c028c",
  1461 => x"050d0402",
  1462 => x"f0050d75",
  1463 => x"881108fe",
  1464 => x"0580cda4",
  1465 => x"082980cd",
  1466 => x"b8081172",
  1467 => x"0880cda8",
  1468 => x"08060579",
  1469 => x"55535454",
  1470 => x"9ec22d02",
  1471 => x"90050d04",
  1472 => x"02f4050d",
  1473 => x"7470882a",
  1474 => x"83fe8006",
  1475 => x"7072982a",
  1476 => x"0772882b",
  1477 => x"87fc8080",
  1478 => x"0673982b",
  1479 => x"81f00a06",
  1480 => x"71730707",
  1481 => x"80c6b80c",
  1482 => x"56515351",
  1483 => x"028c050d",
  1484 => x"0402f805",
  1485 => x"0d028e05",
  1486 => x"80f52d74",
  1487 => x"882b0770",
  1488 => x"83ffff06",
  1489 => x"80c6b80c",
  1490 => x"51028805",
  1491 => x"0d0402f4",
  1492 => x"050d7476",
  1493 => x"78535452",
  1494 => x"80712597",
  1495 => x"38727081",
  1496 => x"055480f5",
  1497 => x"2d727081",
  1498 => x"055481b7",
  1499 => x"2dff1151",
  1500 => x"70eb3880",
  1501 => x"7281b72d",
  1502 => x"028c050d",
  1503 => x"0402e805",
  1504 => x"0d775680",
  1505 => x"70565473",
  1506 => x"7624b638",
  1507 => x"80cdb008",
  1508 => x"742eae38",
  1509 => x"7351a8cf",
  1510 => x"2d80c6b8",
  1511 => x"0880c6b8",
  1512 => x"08098105",
  1513 => x"7080c6b8",
  1514 => x"08079f2a",
  1515 => x"77058117",
  1516 => x"57575353",
  1517 => x"74762489",
  1518 => x"3880cdb0",
  1519 => x"087426d4",
  1520 => x"387280c6",
  1521 => x"b80c0298",
  1522 => x"050d0402",
  1523 => x"f0050d80",
  1524 => x"c6b40816",
  1525 => x"51aefd2d",
  1526 => x"80c6b808",
  1527 => x"802e9f38",
  1528 => x"8b5380c6",
  1529 => x"b8085280",
  1530 => x"cba051ae",
  1531 => x"ce2d80cd",
  1532 => x"dc085473",
  1533 => x"802e8738",
  1534 => x"80cba051",
  1535 => x"732d0290",
  1536 => x"050d0402",
  1537 => x"dc050d80",
  1538 => x"705a5574",
  1539 => x"80c6b408",
  1540 => x"25b43880",
  1541 => x"cdb00875",
  1542 => x"2eac3878",
  1543 => x"51a8cf2d",
  1544 => x"80c6b808",
  1545 => x"09810570",
  1546 => x"80c6b808",
  1547 => x"079f2a76",
  1548 => x"05811b5b",
  1549 => x"56547480",
  1550 => x"c6b40825",
  1551 => x"893880cd",
  1552 => x"b0087926",
  1553 => x"d6388055",
  1554 => x"7880cdb0",
  1555 => x"082781db",
  1556 => x"387851a8",
  1557 => x"cf2d80c6",
  1558 => x"b808802e",
  1559 => x"81ad3880",
  1560 => x"c6b8088b",
  1561 => x"0580f52d",
  1562 => x"70842a70",
  1563 => x"81067710",
  1564 => x"78842b80",
  1565 => x"cba00b80",
  1566 => x"f52d5c5c",
  1567 => x"53515556",
  1568 => x"73802e80",
  1569 => x"cb387416",
  1570 => x"822bb2cf",
  1571 => x"0b80c588",
  1572 => x"120c5477",
  1573 => x"75311080",
  1574 => x"cde01155",
  1575 => x"56907470",
  1576 => x"81055681",
  1577 => x"b72da074",
  1578 => x"81b72d76",
  1579 => x"81ff0681",
  1580 => x"16585473",
  1581 => x"802e8a38",
  1582 => x"9c5380cb",
  1583 => x"a052b1c8",
  1584 => x"048b5380",
  1585 => x"c6b80852",
  1586 => x"80cde216",
  1587 => x"51b28304",
  1588 => x"7416822b",
  1589 => x"afcb0b80",
  1590 => x"c588120c",
  1591 => x"547681ff",
  1592 => x"06811658",
  1593 => x"5473802e",
  1594 => x"8a389c53",
  1595 => x"80cba052",
  1596 => x"b1fa048b",
  1597 => x"5380c6b8",
  1598 => x"08527775",
  1599 => x"311080cd",
  1600 => x"e0055176",
  1601 => x"55aece2d",
  1602 => x"b2a00474",
  1603 => x"90297531",
  1604 => x"701080cd",
  1605 => x"e0055154",
  1606 => x"80c6b808",
  1607 => x"7481b72d",
  1608 => x"81195974",
  1609 => x"8b24a338",
  1610 => x"b0c80474",
  1611 => x"90297531",
  1612 => x"701080cd",
  1613 => x"e0058c77",
  1614 => x"31575154",
  1615 => x"807481b7",
  1616 => x"2d9e14ff",
  1617 => x"16565474",
  1618 => x"f33802a4",
  1619 => x"050d0402",
  1620 => x"fc050d80",
  1621 => x"c6b40813",
  1622 => x"51aefd2d",
  1623 => x"80c6b808",
  1624 => x"802e8938",
  1625 => x"80c6b808",
  1626 => x"51a0a42d",
  1627 => x"800b80c6",
  1628 => x"b40cb083",
  1629 => x"2d918b2d",
  1630 => x"0284050d",
  1631 => x"0402fc05",
  1632 => x"0d725170",
  1633 => x"fd2eb038",
  1634 => x"70fd248a",
  1635 => x"3870fc2e",
  1636 => x"80cc38b3",
  1637 => x"e80470fe",
  1638 => x"2eb73870",
  1639 => x"ff2e0981",
  1640 => x"0680c538",
  1641 => x"80c6b408",
  1642 => x"5170802e",
  1643 => x"bb38ff11",
  1644 => x"80c6b40c",
  1645 => x"b3e80480",
  1646 => x"c6b408f0",
  1647 => x"057080c6",
  1648 => x"b40c5170",
  1649 => x"8025a138",
  1650 => x"800b80c6",
  1651 => x"b40cb3e8",
  1652 => x"0480c6b4",
  1653 => x"08810580",
  1654 => x"c6b40cb3",
  1655 => x"e80480c6",
  1656 => x"b4089005",
  1657 => x"80c6b40c",
  1658 => x"b0832d91",
  1659 => x"8b2d0284",
  1660 => x"050d0402",
  1661 => x"fc050d80",
  1662 => x"0b80c6b4",
  1663 => x"0cb0832d",
  1664 => x"909b2d80",
  1665 => x"c6b80880",
  1666 => x"c6a40c80",
  1667 => x"c5805192",
  1668 => x"ae2d0284",
  1669 => x"050d0471",
  1670 => x"80cddc0c",
  1671 => x"04000000",
  1672 => x"00ffffff",
  1673 => x"ff00ffff",
  1674 => x"ffff00ff",
  1675 => x"ffffff00",
  1676 => x"45786974",
  1677 => x"00000000",
  1678 => x"506f7420",
  1679 => x"33263420",
  1680 => x"4a6f7920",
  1681 => x"32204469",
  1682 => x"73706172",
  1683 => x"6f20322f",
  1684 => x"33000000",
  1685 => x"506f7420",
  1686 => x"33263420",
  1687 => x"5261746f",
  1688 => x"6e000000",
  1689 => x"506f7420",
  1690 => x"33263420",
  1691 => x"50616464",
  1692 => x"6c657320",
  1693 => x"33263400",
  1694 => x"506f7420",
  1695 => x"31263220",
  1696 => x"4a6f7920",
  1697 => x"31204469",
  1698 => x"73706172",
  1699 => x"6f20322f",
  1700 => x"33000000",
  1701 => x"506f7420",
  1702 => x"31263220",
  1703 => x"5261746f",
  1704 => x"6e000000",
  1705 => x"506f7420",
  1706 => x"31263220",
  1707 => x"50616464",
  1708 => x"6c657320",
  1709 => x"31263200",
  1710 => x"50756572",
  1711 => x"746f2055",
  1712 => x"41525400",
  1713 => x"50756572",
  1714 => x"746f204a",
  1715 => x"6f797374",
  1716 => x"69636b73",
  1717 => x"00000000",
  1718 => x"4a6f7973",
  1719 => x"7469636b",
  1720 => x"73204e6f",
  1721 => x"726d616c",
  1722 => x"00000000",
  1723 => x"4a6f7973",
  1724 => x"7469636b",
  1725 => x"7320496e",
  1726 => x"74657263",
  1727 => x"616d6269",
  1728 => x"61646f73",
  1729 => x"00000000",
  1730 => x"4d657a63",
  1731 => x"6c612053",
  1732 => x"74657265",
  1733 => x"6f204e6f",
  1734 => x"00000000",
  1735 => x"4d657a63",
  1736 => x"6c612053",
  1737 => x"74657265",
  1738 => x"6f203235",
  1739 => x"25000000",
  1740 => x"4d657a63",
  1741 => x"6c612053",
  1742 => x"74657265",
  1743 => x"6f203530",
  1744 => x"25000000",
  1745 => x"4d657a63",
  1746 => x"6c612053",
  1747 => x"74657265",
  1748 => x"6f203735",
  1749 => x"25000000",
  1750 => x"45787061",
  1751 => x"6e73696f",
  1752 => x"6e206465",
  1753 => x"20536f6e",
  1754 => x"69646f20",
  1755 => x"4e6f0000",
  1756 => x"45787061",
  1757 => x"6e73696f",
  1758 => x"6e206465",
  1759 => x"20536f6e",
  1760 => x"69646f20",
  1761 => x"4f504c32",
  1762 => x"00000000",
  1763 => x"46696c74",
  1764 => x"726f2064",
  1765 => x"65204175",
  1766 => x"64696f20",
  1767 => x"4f6e0000",
  1768 => x"46696c74",
  1769 => x"726f2064",
  1770 => x"65204175",
  1771 => x"64696f20",
  1772 => x"4f666600",
  1773 => x"53494420",
  1774 => x"44657265",
  1775 => x"63686f20",
  1776 => x"41646472",
  1777 => x"20496775",
  1778 => x"616c0000",
  1779 => x"53494420",
  1780 => x"44657265",
  1781 => x"63686f20",
  1782 => x"41646472",
  1783 => x"20444530",
  1784 => x"30000000",
  1785 => x"53494420",
  1786 => x"44657265",
  1787 => x"63686f20",
  1788 => x"41646472",
  1789 => x"20443432",
  1790 => x"30000000",
  1791 => x"53494420",
  1792 => x"44657265",
  1793 => x"63686f20",
  1794 => x"41646472",
  1795 => x"20443530",
  1796 => x"30000000",
  1797 => x"53494420",
  1798 => x"44657265",
  1799 => x"63686f20",
  1800 => x"41646472",
  1801 => x"20444630",
  1802 => x"30000000",
  1803 => x"53494420",
  1804 => x"44657265",
  1805 => x"63686f20",
  1806 => x"36353831",
  1807 => x"00000000",
  1808 => x"53494420",
  1809 => x"44657265",
  1810 => x"63686f20",
  1811 => x"38353830",
  1812 => x"00000000",
  1813 => x"53494420",
  1814 => x"497a7175",
  1815 => x"69657264",
  1816 => x"6f203635",
  1817 => x"38310000",
  1818 => x"53494420",
  1819 => x"497a7175",
  1820 => x"69657264",
  1821 => x"6f203835",
  1822 => x"38300000",
  1823 => x"5363616e",
  1824 => x"646f7562",
  1825 => x"6c657220",
  1826 => x"4e696e67",
  1827 => x"756e6f00",
  1828 => x"5363616e",
  1829 => x"646f7562",
  1830 => x"6c657220",
  1831 => x"48513278",
  1832 => x"2d333230",
  1833 => x"00000000",
  1834 => x"5363616e",
  1835 => x"646f7562",
  1836 => x"6c657220",
  1837 => x"48513278",
  1838 => x"2d313630",
  1839 => x"00000000",
  1840 => x"5363616e",
  1841 => x"646f7562",
  1842 => x"6c657220",
  1843 => x"43525420",
  1844 => x"32352500",
  1845 => x"5363616e",
  1846 => x"646f7562",
  1847 => x"6c657220",
  1848 => x"43525420",
  1849 => x"35302500",
  1850 => x"5363616e",
  1851 => x"646f7562",
  1852 => x"6c657220",
  1853 => x"43525420",
  1854 => x"37352500",
  1855 => x"466f726d",
  1856 => x"61746f20",
  1857 => x"4f726967",
  1858 => x"696e616c",
  1859 => x"00000000",
  1860 => x"466f726d",
  1861 => x"61746f20",
  1862 => x"50616e74",
  1863 => x"616c6c61",
  1864 => x"20436f6d",
  1865 => x"706c6574",
  1866 => x"61000000",
  1867 => x"466f726d",
  1868 => x"61746f20",
  1869 => x"5b415243",
  1870 => x"315d0000",
  1871 => x"466f726d",
  1872 => x"61746f20",
  1873 => x"5b415243",
  1874 => x"325d0000",
  1875 => x"41737065",
  1876 => x"63746f20",
  1877 => x"4f726967",
  1878 => x"696e616c",
  1879 => x"00000000",
  1880 => x"41737065",
  1881 => x"63746f20",
  1882 => x"416e6368",
  1883 => x"6f000000",
  1884 => x"56696465",
  1885 => x"6f205041",
  1886 => x"4c000000",
  1887 => x"56696465",
  1888 => x"6f204e54",
  1889 => x"53430000",
  1890 => x"2020203d",
  1891 => x"20434f4d",
  1892 => x"4f444f52",
  1893 => x"45202036",
  1894 => x"34203d20",
  1895 => x"20200000",
  1896 => x"20202020",
  1897 => x"20204e65",
  1898 => x"75726f52",
  1899 => x"756c657a",
  1900 => x"20202020",
  1901 => x"20200000",
  1902 => x"20202020",
  1903 => x"20202020",
  1904 => x"20202020",
  1905 => x"20202020",
  1906 => x"20202020",
  1907 => x"20200000",
  1908 => x"52657365",
  1909 => x"74000000",
  1910 => x"52657365",
  1911 => x"74202620",
  1912 => x"536f6c74",
  1913 => x"61722043",
  1914 => x"61727475",
  1915 => x"63686f00",
  1916 => x"56696465",
  1917 => x"6f201000",
  1918 => x"41756469",
  1919 => x"6f201000",
  1920 => x"50756572",
  1921 => x"746f7320",
  1922 => x"10000000",
  1923 => x"53616361",
  1924 => x"72204369",
  1925 => x"6e746100",
  1926 => x"506c6179",
  1927 => x"2f53746f",
  1928 => x"70204369",
  1929 => x"6e746100",
  1930 => x"43617267",
  1931 => x"61722044",
  1932 => x"6973636f",
  1933 => x"2f43696e",
  1934 => x"74612f43",
  1935 => x"61727420",
  1936 => x"10000000",
  1937 => x"44697363",
  1938 => x"6f204772",
  1939 => x"61626162",
  1940 => x"6c650000",
  1941 => x"44697363",
  1942 => x"6f20536f",
  1943 => x"6c6f204c",
  1944 => x"65637475",
  1945 => x"72610000",
  1946 => x"536f6e69",
  1947 => x"646f2043",
  1948 => x"696e7461",
  1949 => x"204f6666",
  1950 => x"00000000",
  1951 => x"536f6e69",
  1952 => x"646f2043",
  1953 => x"696e7461",
  1954 => x"204f6e00",
  1955 => x"4b65726e",
  1956 => x"656c2043",
  1957 => x"61726761",
  1958 => x"626c6500",
  1959 => x"4b65726e",
  1960 => x"656c2043",
  1961 => x"36340000",
  1962 => x"4b65726e",
  1963 => x"656c2043",
  1964 => x"36344753",
  1965 => x"00000000",
  1966 => x"4b65726e",
  1967 => x"656c204a",
  1968 => x"61706f6e",
  1969 => x"65730000",
  1970 => x"43617267",
  1971 => x"61204661",
  1972 => x"6c6c6964",
  1973 => x"61000000",
  1974 => x"4f4b0000",
  1975 => x"16200000",
  1976 => x"14200000",
  1977 => x"15200000",
  1978 => x"53442069",
  1979 => x"6e69742e",
  1980 => x"2e2e0a00",
  1981 => x"53442063",
  1982 => x"61726420",
  1983 => x"72657365",
  1984 => x"74206661",
  1985 => x"696c6564",
  1986 => x"210a0000",
  1987 => x"53444843",
  1988 => x"20657272",
  1989 => x"6f72210a",
  1990 => x"00000000",
  1991 => x"57726974",
  1992 => x"65206661",
  1993 => x"696c6564",
  1994 => x"0a000000",
  1995 => x"52656164",
  1996 => x"20666169",
  1997 => x"6c65640a",
  1998 => x"00000000",
  1999 => x"43617264",
  2000 => x"20696e69",
  2001 => x"74206661",
  2002 => x"696c6564",
  2003 => x"0a000000",
  2004 => x"46415431",
  2005 => x"36202020",
  2006 => x"00000000",
  2007 => x"46415433",
  2008 => x"32202020",
  2009 => x"00000000",
  2010 => x"4e6f2070",
  2011 => x"61727469",
  2012 => x"74696f6e",
  2013 => x"20736967",
  2014 => x"0a000000",
  2015 => x"42616420",
  2016 => x"70617274",
  2017 => x"0a000000",
  2018 => x"4261636b",
  2019 => x"00000000",
  2020 => x"00000002",
  2021 => x"00000003",
  2022 => x"00001ffc",
  2023 => x"00000002",
  2024 => x"00000003",
  2025 => x"00001ff4",
  2026 => x"00000002",
  2027 => x"00000003",
  2028 => x"00001fe8",
  2029 => x"00000003",
  2030 => x"00000003",
  2031 => x"00001fdc",
  2032 => x"00000003",
  2033 => x"00000004",
  2034 => x"00001a30",
  2035 => x"00002128",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00001a38",
  2040 => x"00001a54",
  2041 => x"00001a64",
  2042 => x"00001a78",
  2043 => x"00001a94",
  2044 => x"00001aa4",
  2045 => x"00001ab8",
  2046 => x"00001ac4",
  2047 => x"00001ad8",
  2048 => x"00001aec",
  2049 => x"00000003",
  2050 => x"000020a0",
  2051 => x"00000002",
  2052 => x"00000003",
  2053 => x"00002098",
  2054 => x"00000002",
  2055 => x"00000003",
  2056 => x"00002084",
  2057 => x"00000005",
  2058 => x"00000003",
  2059 => x"0000207c",
  2060 => x"00000002",
  2061 => x"00000003",
  2062 => x"00002074",
  2063 => x"00000002",
  2064 => x"00000003",
  2065 => x"00002064",
  2066 => x"00000004",
  2067 => x"00000004",
  2068 => x"00001a30",
  2069 => x"00002128",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00001b08",
  2074 => x"00001b1c",
  2075 => x"00001b30",
  2076 => x"00001b44",
  2077 => x"00001b58",
  2078 => x"00001b70",
  2079 => x"00001b8c",
  2080 => x"00001ba0",
  2081 => x"00001bb4",
  2082 => x"00001bcc",
  2083 => x"00001be4",
  2084 => x"00001bfc",
  2085 => x"00001c14",
  2086 => x"00001c2c",
  2087 => x"00001c40",
  2088 => x"00001c54",
  2089 => x"00001c68",
  2090 => x"00000003",
  2091 => x"00002120",
  2092 => x"00000002",
  2093 => x"00000003",
  2094 => x"00002118",
  2095 => x"00000002",
  2096 => x"00000003",
  2097 => x"00002108",
  2098 => x"00000004",
  2099 => x"00000003",
  2100 => x"000020f0",
  2101 => x"00000006",
  2102 => x"00000004",
  2103 => x"00001a30",
  2104 => x"00002128",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00001c7c",
  2109 => x"00001c90",
  2110 => x"00001ca8",
  2111 => x"00001cc0",
  2112 => x"00001cd4",
  2113 => x"00001ce8",
  2114 => x"00001cfc",
  2115 => x"00001d10",
  2116 => x"00001d2c",
  2117 => x"00001d3c",
  2118 => x"00001d4c",
  2119 => x"00001d60",
  2120 => x"00001d70",
  2121 => x"00001d7c",
  2122 => x"00000002",
  2123 => x"00001d88",
  2124 => x"00000000",
  2125 => x"00000002",
  2126 => x"00001da0",
  2127 => x"00000000",
  2128 => x"00000002",
  2129 => x"00001db8",
  2130 => x"00000000",
  2131 => x"00000002",
  2132 => x"00001dd0",
  2133 => x"00000371",
  2134 => x"00000002",
  2135 => x"00001dd8",
  2136 => x"00000388",
  2137 => x"00000004",
  2138 => x"00001df0",
  2139 => x"000020a8",
  2140 => x"00000004",
  2141 => x"00001df8",
  2142 => x"00002004",
  2143 => x"00000004",
  2144 => x"00001e00",
  2145 => x"00001f94",
  2146 => x"00000003",
  2147 => x"000021f8",
  2148 => x"00000004",
  2149 => x"00000003",
  2150 => x"000021f0",
  2151 => x"00000002",
  2152 => x"00000003",
  2153 => x"000021e8",
  2154 => x"00000002",
  2155 => x"00000002",
  2156 => x"00001e0c",
  2157 => x"000003b8",
  2158 => x"00000002",
  2159 => x"00001e18",
  2160 => x"000003a0",
  2161 => x"00000002",
  2162 => x"00001e28",
  2163 => x"000019f3",
  2164 => x"00000002",
  2165 => x"00001a30",
  2166 => x"00000824",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00001e44",
  2171 => x"00001e54",
  2172 => x"00001e68",
  2173 => x"00001e7c",
  2174 => x"00001e8c",
  2175 => x"00001e9c",
  2176 => x"00001ea8",
  2177 => x"00001eb8",
  2178 => x"00000004",
  2179 => x"00001ec8",
  2180 => x"00002208",
  2181 => x"00000004",
  2182 => x"00001ed8",
  2183 => x"00002128",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"00000002",
  2209 => x"000026e0",
  2210 => x"000017cb",
  2211 => x"00000002",
  2212 => x"000026fe",
  2213 => x"000017cb",
  2214 => x"00000002",
  2215 => x"0000271c",
  2216 => x"000017cb",
  2217 => x"00000002",
  2218 => x"0000273a",
  2219 => x"000017cb",
  2220 => x"00000002",
  2221 => x"00002758",
  2222 => x"000017cb",
  2223 => x"00000002",
  2224 => x"00002776",
  2225 => x"000017cb",
  2226 => x"00000002",
  2227 => x"00002794",
  2228 => x"000017cb",
  2229 => x"00000002",
  2230 => x"000027b2",
  2231 => x"000017cb",
  2232 => x"00000002",
  2233 => x"000027d0",
  2234 => x"000017cb",
  2235 => x"00000002",
  2236 => x"000027ee",
  2237 => x"000017cb",
  2238 => x"00000002",
  2239 => x"0000280c",
  2240 => x"000017cb",
  2241 => x"00000002",
  2242 => x"0000282a",
  2243 => x"000017cb",
  2244 => x"00000002",
  2245 => x"00002848",
  2246 => x"000017cb",
  2247 => x"00000004",
  2248 => x"00001f88",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"0000197d",
  2253 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

